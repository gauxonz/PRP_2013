************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA85
* BEGIN OPAMP MACROMODEL PA93
* NOTE THAT IQ PIN IS NOT MODELED
* PINOUT ORDER +IN -IN CL OUT +V -V COMP COMP
*                1   2  3  33  4  5   6    7
.SUBCKT PA93 1 2 3 33 4 5 6 7
J1 10 1 8 JI1
J2 11 36 9 JI2
R3 12 8 5.17E+02
R4 12 9 5.17E+02
I2 12 5 7.2E-04
C1 12 5 4.32E-13
R5 12 5 9.72E+07
C7 9 41 3.08E-10
RZ1 12 40 5.17E+01
C8 8 40 3.08E-10
RZ2 12 41 5.17E+01
R1 4 10 5.42E+02
R2 4 11 5.42E+02
C2 10 11 5.88E-11
I1 4 5 -6.91E-03
G1 6 15 11 10 1.85E-03
G2 37 15 12 15 1.00E-04
LCM 37 38 1.0E-06
RCM 15 38 1.0
ECA 2 36 37 15 1.0
R6 6 15 1.00E+05
D1 6 34 DD
D7 34 15 DD
D2 35 6 DD
D8 15 35 DD
C3 6 7 4.70E-12
G3 15 7 15 6 3.42E-01
R7 7 15 1E3
D3 7 16 DD
V1 18 16 6.20E+00
D4 17 7 DD
V2 17 19 6.20E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 42 50
C4 42 15 2.80E-11
R11 20 42 50
C5 20 15 6.37E-10
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 333
R10 28 3 333
I3 18 21 1.64E-02
I4 22 19 1.64E-02
R15 29 3 3.43E-01
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=1.57E-13 RS=1.90E-02)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL JI1 NJF (BETA=4.00E-02 IS=3E-16 VTO=-1 KF=7.0E-18)
.MODEL JI2 NJF (BETA=4.00E-02 IS=3E-16 VTO=-1.0020 KF=7.0E-18)
.MODEL QOP PNP (BF=9.60E+02 IS=1E-14)
.MODEL QON NPN (BF=9.60E+02 IS=1E-14)
.MODEL QLN NPN (BF=200 IS=6E-13)
.MODEL QLP PNP (BF=200 IS=6E-13)
* END OF OPAMP MACROMODEL
.ENDS
*************
