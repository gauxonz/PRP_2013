* Readme.txt
*       THESE MODELS ARE PROVIDED AS IS WITH NO WARRANTY STATED
*	OR IMPLIED. NIETHER APEX MICROTECHNOLOGY NOR ANALOG AND
*       RF MODELS SHALL BE HELD LIABLE FOR ANY DAMAGES RELATING
*	TO THE USE OF THESE MODELS.
*
*
*       MOST APEX LINEAR SPICE MODES ARE COMPATIBLE WITH
*       BOTH PSPICE AND BERKELEY DERIVED SIMULATORS.  THEY ARE
*       PROVIDED IN BOTH INDIVIDUAL FILES AND A TOTAL FILE FOR
*       USER CONVENIENCE.  THERE IS NO DIFFERENCE BETWEEN MODELS
*       OF THE TWO GROUPS.  THIS FILE APPEARS AT THE TOP OF
*       THE TOTAL FILE.  IT IS NOT REPEATED IN THE INDIVIDUAL
*       FILES, BUT APPLIES TO EACH.
*
*       THE PA69, PA78, PA86, PA240, PA241 AND PA243 MODELS CONTAIN  
*       RESISTORS WITH TEMPERATURE COEFFICIENTS THAT REQUIRE DIFFERENT 
*       SYNTAX FOR PSPICE AND BERKELEY DERIVED SIMULATORS.  THESE
*       MODELS ARE CONTAINED IN SEPARATE .ZIP FILES. BE AWARE THAT
*       THE MODELS INSIDE THESE TWO FILES HAVE IDENTICAL NAMES.  OTHER
*       MODELS ARE COMPATIBLE WITH EITHER TYPE SIMULATOR.     
*
************
*   FEATURES OF THE APEX OP AMP MACROMODELS FOR SPICE
*
*	THE APEX MACROMODELS ELIMINATE MANY OF THE CONVERGENCE
*	AND TIMESTEP PROBLEMS OF AN EXACT MODEL WHILE EXECUTING
*	MANY TIMES FASTER DURING SIMULATION. IN SOME CIRCUITS
*	DC CONVERGENCE WILL REQUIRE THAT THE OP AMP OUTPUT BE
*	NODESET NEAR ITS OPERATING POINT. USING FEEDBACK FROM
*	CUSTOMERS, WE HAVE ATTEMPTED TO OFFER THE BEST PRACTICAL
*	TRADEOFF OF FEATURES, REALISM, COMPLEXITY, EASE OF USE,
*	COMPATIBILITY WITH COMMONLY AVAILABLE SPICE SIMULATORS,
*	AND SIMULATION RUN TIME IN THESE MACROMODELS. SOME SIM-
*	ULATORS MAY REQUIRE MINOR SYNTAX EDITING.  MODELS 
*       FUNCTION UNDER SPICE 2G.6 OR 3X.X
*
*   CHARACTERISTICS MODELED :
*
*	 1 PROPER OPEN LOOP GAIN AND PHASE
*	 2 PROPER UNSYMMETRICAL OUTPUT VOLTAGE SWING
*	 3 PROPER SMALL SIGNAL OPEN LOOP OUTPUT IMPEDANCE (SSZO)
*	 4 PROPER OUTPUT VOLTAGE SWING DROOP WITH OUTPUT CURRENT
*	   (LSZO)
*	 5 PROPER TRANSITION OF OUTPUT IMPEDANCE FROM
*	   SSZO TO LSZO AS OUTPUT CURRENT RISES
*	 6 PROPER QUIESCENT CURRENT THROUGH SUPPLY PINS
*	 7 OUTPUT CURRENT FLOW THROUGH THE SUPPLY PINS
*	 8 PROPER OUTPUT CURRENT LIMIT CHARACTERISTICS
*	   VERSUS TEMPERATURE
*	 9 REALISTIC SATURATION RECOVERY TIME
*	10 REALISTIC COMPENSATION
*	11 REALISTIC UNSYMMETRICAL SLEW RATE
*	12 INPUT COMMON MODE REJECTION
*	13 BIPOLAR, JFET, OR MOSFET INPUT STAGE DEPENDING
*	   ON THE REAL PART
*	14 OUTPUT TO SUPPLY CLAMPING DIODES DEPENDING ON
*	   THE REAL PART AND INTERNAL MOSFET CLAMP DIODES,
*	   IF THE REAL PART HAS MOSFET OUTPUT DEVICES
*	15 INPUT OFFSET VOLTAGE
*	16 INPUT BIAS CURRENT AND OFFSET IF BIPOLAR FRONT END
*	17 USE NO INTERNAL POLYNOMIAL SOURCES
*	18 OPERATION OVER TEMPERATURE
*	19 NO REQUIREMENT FOR A GROUND REFERENCE
*	20 PROPER MAXIMUM OUTPUT CURRENT IF CURRENT LIMIT
*	   RESISTOR(S) ARE SMALLER THAN MINIMUM ALLOWED
*	21 IMPROVED CMRR VS FREQUENCY IS MODELED IN THE
*	   PA90, PA91, PA92, PA93 ONLY
*
*   CHARACTERISTICS NOT MODELED :
*
*	 1 INPUT BIAS CURRENT FOR JFET AND MOSFET INPUT TYPES
*	 2 INPUT AND OUTPUT CAPACITANCE
*	 3 POWER SUPPLY REJECTION
*	 4 EXACT FREQUENCY PROFILE OF CMRR
*	 5 EXACT HARMONIC DISTORTION
*	 6 EXACT INPUT COMMON MODE VOLTAGE RANGE
*	 7 MIN OR MAX POWER SUPPLY VOLTAGE FAILURE
*	 8 OFFSET BALANCE PINS NOT INCLUDED
*	 9 INPUT VOLTAGE AND CURRENT NOISE
*	10 IQ PIN NOT MODELED
*
*
*   MACROMODELS INCLUDED IN THIS FILE:
*	MA01, MP38, MP39, PA01, PA02, PA03, PA04, PA05, PA07, 
*	PA08, PA09, PA10, PA12, PA13, PA140, PA141, PA142, PA144,
*	PA15, PA16, PA162,PA19, PA21, PA25, PA26, PA33, PA34, PA35AMP,
*	PA35BUF, PA37, PA40, PA41, PA42, PA44, PA50, PA51, PA52,
*	PA60, PA61, PA62, PA73, PA74, PA75AMP, PA75BUF, PA76, PA81,
*	PA83, PA84, PA85, PA88, PA89, PA90, PA91, PA92, PA93, PA94,
*	PA95, PA97, PA98, PA240, PA241, PB50, PB51, PB51A, PB58, PB58A
*
*   NOTE: WHEN USING PA26, PA34 OR PA37 WITHOUT VBOOST OR ISENSE
*       FEATURES, THE PA25 HAVING 2 LESS PINS WILL WORK.
* 
**************
*
*   FEATURES OF THE APEX OP AMP ENHANCED MODELS FOR SPICE
*	THE APEX ENHANCED MODELS ARE MOSTLY COMPONENT BASED TO
*	ADD ACCURACY AND FEATURES.  GREAT CARE WAS TAKEN TO AVOID
*	CONVERGENCE AND TIMESTEP PROBLEMS OR EXCESSIVE RUN TIMES. 
*	IN SOME CIRCUITS DC CONVERGENCE WILL REQUIRE THAT THE OP 
*	AMP OUTPUT BE NODESET NEAR ITS OPERATING POINT.  SOME SIM-
*	ULATORS MAY REQUIRE MINOR SYNTAX EDITING.  MODELS 
*       FUNCTION UNDER SPICE 3X.X
*
*
*   CHARACTERISTICS MODELED :
*
*	 1 ALL PARAMETERS LISTED FOR MACROMODELS
*	 2 INPUT AND OUTPUT CAPACITANCE
*	 3 POWER SUPPLY REJECTION
*	 4 FREQUENCY PROFILE OF CMRR
*	 5 HARMONIC DISTORTION
*	 6 INPUT COMMON MODE VOLTAGE RANGE
*	 7 MIN OR MAX POWER SUPPLY VOLTAGE FAILURE
*	 8 SHUTDOWN IF APPLICABLE
*	 9 IQ PIN IF APPLICABLE
*
*   CHARACTERISTICS NOT MODELED :
*
*	 1 INPUT VOLTAGE AND CURRENT NOISE
*
*   ENHANCED MODELS INCLUDED IN THIS FILE:
*
*        MP38, MP39, MP108, MP111,MP230, MP240, PA69, PA78, PA79, PA86
*
*************
*
*	FOR OTHER SPICE MODELS EMAIL ANALOG AND RF MODELS,
*       WKSANDS@EARTHLINK.NET.
*
*************************
*SYM=PA85
* BEGIN OPAMP MACROMODEL MA01
* PINOUT ORDER +IN -IN CL OUT +V -V COMP COMP
*                1   2  3  33  4  5   6    7
.SUBCKT MA01 1 2 3 33 4 5 6 7
M1 10 1 8 8 MI1
M2 11 2 9 9 MI2
R3 12 8 2.95E+03
R4 12 9 2.95E+03
I2 12 5 2.90E-04
C1 12 5 7.78E-13
R5 12 5 1.38E+07
R1 4 10 3.20E+03
R2 4 11 3.20E+03
C2 10 11 1.66E-11
I1 4 5 -8.81E-05
G1 6 15 11 10 3.13E-04
G2 6 15 12 15 5.56E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 5.00E-12
G3 15 7 15 6 5.69E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 3.20E+00
D4 17 7 DD
V2 17 19 6.70E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 9.35E-11
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
M3 25 27 33 33 MLN
M4 26 28 33 33 MLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 1.20E-03
I4 22 19 1.20E-03
R15 29 3 7.50E+01
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=8.40E-16 RS=3.57E+00)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MI1 NMOS (KP=4.00E-03 IS=3E-16 VTO=1)
.MODEL MI2 NMOS (KP=4.00E-03 IS=3E-16 VTO=0.9850)
.MODEL MLN NMOS (KP=5.00E-03 IS=3E-16 VTO=2.5)
.MODEL MLP PMOS (KP=5.00E-03 IS=3E-16 VTO=-2.5)
.MODEL QOP PNP (BF=7.01E+01 IS=1E-14)
.MODEL QON NPN (BF=7.01E+01 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
*************
* REVISION 1 9-OCT-2006
* BEGIN MODEL MP108
* PINOUT ORDER +IN -IN +ILIM -ILIM OUT +VB -VB
*               1   2    5     4    3   6   7
*              COMP COMP +VS -VS
*                8    9   10  11
* NOTE THAT UPPER AND LOWER FETS ARE BROUGHT
* TO THE OUTPUT ON ONE PIN IN THE MODEL
.SUBCKT MP108 1 2 5 4 3 6 7 8 9 10 11
X1 10 12 13 IRF640NS
X7 11 14 15 IRF9640
R77 16 6 15
C1 6 17 470E-12
R83 18 12 10
R85 19 14 10
R86 9 20 100
R93 7 21 350
R94 7 22 113
Q12 8 16 6 Q907
D6 8 6 C8V2
E2 23 24 6 7 -30E-6
D8 25 0 DD
I1 0 25 1E-3
V16 25 26 0.7
E3 27 0 26 0 -571
R98 0 26 1E6
R99 0 27 1E6
E4 28 18 29 0 -1E-7
E5 30 19 29 0 1E-7
V17 27 29 27
R100 0 29 1E6
D9 23 31 DZ
D10 32 33 C5V6
J2 32 34 35 N912
J3 8 36 37 N912
R101 38 35 30
R102 38 37 30
Q13 33 39 40 Q907B
Q14 8 33 41 Q907B
R103 40 6 82.5
R104 41 6 82.5
J4 8 32 8 N912
R105 32 33 1E5
D11 40 6 C8V2
V18 36 42 -5.75E-3
R106 33 39 70
R109 17 16 120
Q15 43 44 4 Q222
Q16 45 44 4 Q908
R110 44 5 100
R116 2 34 10
R117 1 46 10
C4 6 47 470E-12
C5 47 7 470E-12
E99 48 49 50 0 0.15
R118 50 51 1E6
R119 0 50 100
C25 51 50 1E-12
E100 51 0 6 0 1
R120 49 48 1E9
E101 49 52 53 0 -0.15
R121 53 54 1E6
R122 0 53 100
C26 54 53 20E-12
E102 54 0 7 0 1
R123 52 49 1E9
E103 52 55 56 0 -0.14
R124 56 57 1E6
R125 0 56 100
C27 57 56 20E-12
E104 57 0 58 0 1
R126 55 52 1E9
E105 55 46 59 60 4
D17 59 0 DVN
I7 0 59 100E-6
D18 60 0 DVN
I8 0 60 100E-6
R127 46 55 1E9
E106 61 0 48 0 1
E107 62 0 34 0 1
R128 58 61 1E3
R129 58 62 1E3
R130 7 6 12E3
E108 42 48 29 0 50E-6
R131 48 42 1E9
C28 34 0 2E-12
C29 48 0 2E-12
I9 6 7 -2E-3
R133 24 23 1E9
X10 63 7 22 D560
X11 38 7 21 D560
X12 20 8 17 P450
R134 0 47 1
R145 13 3 0.005
R148 15 3 0.03
Q17 6 20 64 F458
Q18 7 31 65 F558
Q19 66 66 20 F558
Q20 66 66 31 F458
Q21 6 24 67 F458
Q22 7 63 68 F558
Q23 69 69 24 F558
Q24 69 69 63 F458
R149 28 64 6
R150 65 28 6
R151 30 67 6
R152 68 30 6
C31 31 24 2200E-12
C32 8 9 4.6E-12
D19 20 43 D48
D20 45 24 D48
C33 44 45 4700E-12
C34 43 44 4700E-12
R155 0 19 1E12
R156 0 18 1E12
.MODEL D48 D RS=10 IS=1E-15 CJO=1E-12 TT=1N
.MODEL F458  NPN BF=210 IKF=0.5 VAF=1050
+XTB=1.4 ISE=2.1E-14
+ISC=6.42E-12  RB=0.5 RE=0.224 RC=0.134 CJC=12.75E-12
+MJC=0.3966 VJC=0.4332 CJE=183E-12 TF=2.49E-9
.MODEL F558 PNP BF=200 IKF=0.5 VAF=349
+ISE=3.35E-14  ISC=9.42E-12
+ RB=0.133 RE=0.5725 RC=0.748 CJC=26.4E-12 MJC=0.5932 
+VJC=0.9135 CJE=165E-12 TF=1.7E-9
.MODEL DVN D KF=5E-16
.MODEL DD D
.MODEL MSD PMOS KP=0.05 VTO=-2
.MODEL Q222 NPN IS=2E-13
.MODEL Q908 PNP IS=1E-13
.MODEL DZ D BV=6.135 IBV=0.001 RS=5
.MODEL N912 NJF VTO=-3 BETA=3.2E-3 RS=12 RD=50
+ IS=1E-18 LAMBDA=3E-4 CGS=10E-12 CGD=0.5E-12
.MODEL C5V6 D IS=1E-15 RS=5 N=1 BV=5.6 IBV=1E-4
.MODEL C8V2 D IS=1E-15 RS=5 N=1 BV=8.2 IBV=1E-4
.MODEL Q907 PNP IS=1.1E-13 BF=150 BR=6 NF=1.2
+ RC=1 IKF=0.1 VAF=90 XTB=1.5 NE=1.8 ISE=1.5E-13
+ CJE=20E-12 VJE=0.8 MJE=1.2 CJC=15E-12 VJC=0.57
+ MJC=0.3 TF=0.5E-9 TR=35E-9
.MODEL Q907B PNP IS=1.1E-13 BF=150 BR=6 NF=1.2
+ RC=1 IKF=0.1 VAF=900 XTB=1.5 NE=1.8 ISE=1.5E-13
+ CJE=20E-12 VJE=0.8 MJE=1.2 CJC=15E-12 VJC=0.57
+ MJC=0.3 TF=0.5E-9 TR=35E-9
.ENDS MP108
.SUBCKT D560 10 20 30
M1 10 20 30 30 DMOS L=1U W=1U
CGS 20 30 43E-12
.MODEL DMOS NMOS LEVEL=3 VMAX=9E5 THETA=6E-3 ETA=2E-4
+ VTO=-2.5 KP=0.07 RS=2 RD=19)
.ENDS
.SUBCKT P450 10 20 30
M1 10 20 30 30 DMOS L=1U W=1U
RDS 10 30 1E6
CGS 20 30 85E-12
CDG 10 20 20E-12
.MODEL DMOS PMOS LEVEL=3 VMAX=9E5 THETA=60E-3 ETA=2E-3
+ VTO=-2 KP=0.05 RS=3 RD=10)
.ENDS
.SUBCKT irf640ns 1 2 3
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on Feb 14, 02
* MODEL FORMAT: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
.MODEL MM NMOS LEVEL=1 IS=1e-32
+VTO=4.12428 LAMBDA=0.00426564 KP=7.74523
+CGSO=1.06e-05 CGDO=1e-10
RS 8 3 1e-05
D1 3 1 MD
.MODEL MD D IS=4.09854e-11 RS=0.00724292 N=1.17043 BV=200
+IBV=0.00025 EG=1.2 XTI=4 TT=0
+CJO=8e-10 VJ=1.41926 M=0.676432 FC=0.5
RDS 3 1 1e+06
RD 9 1 0.1
RG 2 7 1.35527
D2 4 5 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=1.5322e-09 VJ=1.34184 M=0.9 FC=1e-08
D3 0 5 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=3e-15 N=0.693912 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 2.19598e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=3e-15 N=0.693912
.ENDS
.SUBCKT irf9640 1 2 3
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on May 21, 96
* Model format: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
* Default values used in MM:
* The voltage-dependent capacitances are
* not included. Other default values are:
*   RS=0 RD=0 LD=0 CBD=0 CBS=0 CGBO=0
.MODEL MM PMOS LEVEL=1 IS=1e-32
+VTO=-3.8062 LAMBDA=0.0228396 KP=10.7224
+CGSO=1.09465e-05 CGDO=1e-11
RS 8 3 0.101556
D1 1 3 MD
.MODEL MD D IS=1e-17 RS=0.185714 N=1.5 BV=200
+IBV=0.00025 EG=1.2 XTI=4 TT=1e-07
+CJO=1.22255e-09 VJ=2.42988 M=0.605683 FC=0.493595
RDS 3 1 2e+06
RD 9 1 0.261579
RG 2 7 6.81119
D2 5 4 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=8.6947e-10 VJ=2.34088 M=0.9 FC=1e-08
D3 5 0 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=3e-15 N=0.402798 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 1.8148e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 6 0 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=3e-15 N=0.402798
.ENDS
* END MODEL MP108
*************
* REVISION 1 9-OCT-2006
* BEGIN MODEL MP111
* PINOUT ORDER +IN -IN +ILIM -ILIM OUT +VB -VB
*               1   2    5     4    3   6   7
*              COMP COMP +VS -VS
*                8    9   10  11
* NOTE THAT UPPER AND LOWER FETS ARE BROUGHT
* TO THE OUTPUT ON ONE PIN IN THE MODEL
.SUBCKT MP111 1 2 5 4 3 6 7 8 9 10 11
X1 10 12 13 IRF3710S
X7 11 14 15 IRF5210S
R77 16 6 15
C1 6 17 470E-12
R83 18 12 10
R85 19 14 10
R86 9 20 100
R93 7 21 350
R94 7 22 113
Q12 8 16 6 Q907
D6 8 6 C8V2
E2 23 24 6 7 -30E-6
D8 25 0 DD
I1 0 25 1E-3
V16 25 26 0.7
E3 27 0 26 0 -571
R98 0 26 1E6
R99 0 27 1E6
E4 28 18 29 0 -135E-6
E5 30 19 29 0 135E-6
V17 27 29 27
R100 0 29 1E6
D9 23 31 DZ
D10 32 33 C5V6
J2 32 34 35 N912
J3 8 36 37 N912
R101 38 35 30
R102 38 37 30
Q13 33 39 40 Q907B
Q14 8 33 41 Q907B
R103 40 6 82.5
R104 41 6 82.5
J4 8 32 8 N912
R105 32 33 1E5
D11 40 6 C8V2
V18 36 42 -5.25E-3
R106 33 39 70
R109 17 16 120
Q15 43 44 4 Q222
Q16 45 44 4 Q908
R110 44 5 100
R116 2 34 10
R117 1 46 10
C4 6 47 470E-12
C5 47 7 470E-12
E99 48 49 50 0 0.15
R118 50 51 1E6
R119 0 50 100
C25 51 50 1E-12
E100 51 0 6 0 1
R120 49 48 1E9
E101 49 52 53 0 -0.15
R121 53 54 1E6
R122 0 53 100
C26 54 53 20E-12
E102 54 0 7 0 1
R123 52 49 1E9
E103 52 55 56 0 -0.14
R124 56 57 1E6
R125 0 56 100
C27 57 56 20E-12
E104 57 0 58 0 1
R126 55 52 1E9
E105 55 46 59 60 4
D17 59 0 DVN
I7 0 59 100E-6
D18 60 0 DVN
I8 0 60 100E-6
R127 46 55 1E9
E106 61 0 48 0 1
E107 62 0 34 0 1
R128 58 61 1E3
R129 58 62 1E3
R130 7 6 3.5E3
E108 42 48 29 0 50E-6
R131 48 42 1E9
C28 34 0 2E-12
C29 48 0 2E-12
I9 6 7 -7E-3
R133 24 23 1E9
X10 63 7 22 D560
X11 38 7 21 D560
X12 20 8 17 P450B
R134 0 47 1
R145 13 3 0.043
R148 15 3 0.001
Q17 6 20 64 F458
Q18 7 31 65 F558
Q19 66 66 20 F558
Q20 66 66 31 F458
Q21 6 24 67 F458
Q22 7 63 68 F558
Q23 69 69 24 F558
Q24 69 69 63 F458
R149 28 64 2
R150 65 28 2
R151 30 67 2
R152 68 30 2
C31 31 24 2200E-12
C32 8 9 3E-12
D19 20 43 D48
D20 45 24 D48
C34 43 44 4700E-12
C35 44 45 4700E-12
R158 0 18 1E12
R159 0 19 1E12
.MODEL D48 D RS=10 IS=1E-15 CJO=1E-12 TT=1N
.MODEL F458  NPN BF=210 IKF=0.5 VAF=1050
+XTB=1.4 ISE=2.1E-14
+ISC=6.42E-12  RB=0.5 RE=0.224 RC=0.134 CJC=12.75E-12
+MJC=0.3966 VJC=0.4332 CJE=183E-12 TF=2.49E-9
.MODEL F558 PNP BF=200 IKF=0.5 VAF=349
+ISE=3.35E-14  ISC=9.42E-12
+ RB=0.133 RE=0.5725 RC=0.748 CJC=26.4E-12 MJC=0.5932 
+VJC=0.9135 CJE=165E-12 TF=1.7E-9
.MODEL DVN D KF=5E-16
.MODEL DD D
.MODEL MSD PMOS KP=0.05 VTO=-2
.MODEL Q222 NPN IS=2E-13
.MODEL Q908 PNP IS=1E-13
.MODEL DZ D BV=5.86 IBV=0.001 RS=5
.MODEL N912 NJF VTO=-3 BETA=3.2E-3 RS=12 RD=50
+ IS=1E-18 LAMBDA=3E-4 CGS=10E-12 CGD=0.5E-12
.MODEL C5V6 D IS=1E-15 RS=5 N=1 BV=5.6 IBV=1E-4
.MODEL C8V2 D IS=1E-15 RS=5 N=1 BV=8.2 IBV=1E-4
.MODEL Q907 PNP IS=1.1E-13 BF=150 BR=6 NF=1.2
+ RC=1 IKF=0.1 VAF=90 XTB=1.5 NE=1.8 ISE=1.5E-13
+ CJE=20E-12 VJE=0.8 MJE=1.2 CJC=15E-12 VJC=0.57
+ MJC=0.3 TF=0.5E-9 TR=35E-9
.MODEL Q907B PNP IS=1.1E-13 BF=150 BR=6 NF=1.2
+ RC=1 IKF=0.1 VAF=900 XTB=1.5 NE=1.8 ISE=1.5E-13
+ CJE=20E-12 VJE=0.8 MJE=1.2 CJC=15E-12 VJC=0.57
+ MJC=0.3 TF=0.5E-9 TR=35E-9
.ENDS MP111
.SUBCKT D560 10 20 30
M1 10 20 30 30 DMOS L=1U W=1U
CGS 20 30 43E-12
.MODEL DMOS NMOS LEVEL=3 VMAX=9E5 THETA=6E-3 ETA=2E-4
+ VTO=-2.5 KP=0.07 RS=2 RD=19
.ENDS
.SUBCKT P450B 10 20 30
M1 10 20 30 30 DMOS L=1U W=1U
RDS 10 30 1E6
CGS 20 30 85E-12
CDG 10 20 10E-12
.MODEL DMOS PMOS LEVEL=3 VMAX=9E5 THETA=60E-3 ETA=2E-3
+ VTO=-2 KP=0.05 RS=3 RD=10)
.ENDS
.SUBCKT irf3710s 1 2 3
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on Apr 24, 96
* Model format: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
* Default values used in MM:
* The voltage-dependent capacitances are
* not included. Other default values are:
*   RS=0 RD=0 LD=0 CBD=0 CBS=0 CGBO=0
.MODEL MM NMOS LEVEL=1 IS=1e-32
+VTO=3.73708 LAMBDA=0 KP=46.8579
+CGSO=2.80329e-05 CGDO=1.13722e-06
RS 8 3 0.0113627
D1 3 1 MD
.MODEL MD D IS=9.43288e-12 RS=0.00528331 N=1.07071 BV=100
+IBV=0.00025 EG=1 XTI=3.04957 TT=1e-07
+CJO=1.84661e-09 VJ=0.520811 M=0.45842 FC=0.1
RDS 3 1 4e+06
RD 9 1 0.00538705
RG 2 7 3.87439
D2 4 5 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=4.17518e-09 VJ=0.5 M=0.749785 FC=1e-08
D3 0 5 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=3e-15 N=0.40022 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 6.93446e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=1e-10 N=0.40022
.ENDS
.SUBCKT irf5210s 1 2 3
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on Apr 23, 96
* Model format: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
* Default values used in MM:
* The voltage-dependent capacitances are
* not included. Other default values are:
*   RS=0 RD=0 LD=0 CBD=0 CBS=0 CGBO=0
.MODEL MM PMOS LEVEL=1 IS=1e-32
+VTO=-3.79917 LAMBDA=0.00220079 KP=12.9564
+CGSO=2.34655e-05 CGDO=1e-11
RS 8 3 0.0218795
D1 1 3 MD
.MODEL MD D IS=2.06405e-13 RS=0.00826096 N=0.960301 BV=100
+IBV=0.00025 EG=1 XTI=3.14871 TT=1e-07
+CJO=1.88397e-09 VJ=1.14128 M=0.533786 FC=0.1
RDS 3 1 4e+06
RD 9 1 0.014128
RG 2 7 7.71191
D2 5 4 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=4.75211e-09 VJ=1.32261 M=0.798237 FC=1e-08
D3 5 0 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=3e-15 N=0.40011 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 6.15698e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 6 0 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=1e-10 N=0.40011
.ENDS
* END MODEL MP111
*************
* REVISION 1 29-NOV-2005
* BEGIN MODEL MP230
* PINOUT ORDER +IN -IN +VB -VB GND CC1 CC2 IQ LSD HSD
*               41  42  1   38  2   6   4   5  7   8
*              +VS RS1 RS2 +ILIM -ILIM RS3 RS4 -VS
*               12  9   15   36    35   24  30  21
*
.SUBCKT MP230 41 42 1 38 2 6 4 5 7 8 12 9 15 36 35 24 30 21
X1 12 43 44 IRF540NS
X7 21 45 46 IRF9540N
R77 47 1 20
C1 1 48 470E-12
X8 12 49 50 IRF540NS
X9 21 51 52 IRF9540N
R82 53 49 10
R83 53 43 10
R84 54 51 10
R85 54 45 10
R86 6 55 100
R93 38 56 425
R94 38 57 157
Q12 4 47 1 Q907
D6 4 1 C8V2
E2 58 5 1 38 -5E-6
D8 59 0 DD
I1 0 59 1E-3
V16 59 60 0.7
E3 61 0 60 0 -571
R98 0 60 1E6
R99 0 61 1E6
E4 53 55 0 62 1.135E-3
E5 54 5 62 0 1.135E-3
V17 61 62 27
R100 0 62 1E6
D9 58 55 DZ
D10 63 64 C5V6
J2 63 65 66 N912
J3 4 67 68 N912
R101 69 66 30
R102 69 68 30
Q13 64 70 71 Q907
Q14 4 64 72 Q907
R103 71 1 100
R104 72 1 100
J4 4 63 4 N912
R105 63 64 1E5
D11 71 1 C8V2
V18 67 73 -0.5E-3
R106 64 70 160
C3 53 54 0.01E-6
R109 48 47 75
Q15 74 75 35 Q222
Q16 76 75 35 Q908
R110 75 36 100
Q17 76 52 77 Q908
R111 77 78 130
R112 77 79 5.1
Q18 74 78 79 Q222
R113 80 1 7000
Q20 80 8 81 Q222
R115 7 81 2700
D15 53 74 C5V6
D16 76 54 C5V6
R116 42 65 10
R117 41 82 10
C4 1 2 470E-12
C5 2 38 470E-12
E99 83 84 85 0 0.15
R118 85 86 1E6
R119 0 85 100
C25 86 85 1E-12
E100 86 0 1 0 1
R120 84 83 1E9
E101 84 87 88 0 0.15
R121 88 89 1E6
R122 0 88 100
C26 89 88 20E-12
E102 89 0 38 0 1
R123 87 84 1E9
E103 87 90 91 0 -0.15
R124 91 92 1E6
R125 0 91 100
C27 92 91 20E-12
E104 92 0 93 0 1
R126 90 87 1E9
E105 90 82 94 95 4
D17 94 0 DVN
I7 0 94 100E-6
D18 95 0 DVN
I8 0 95 100E-6
R127 82 90 1E9
E106 96 0 83 0 1
E107 97 0 65 0 1
R128 93 96 1E3
R129 93 97 1E3
R130 38 1 50E3
E108 73 83 62 0 5E-6
R131 83 73 1E9
C28 65 0 2E-12
C29 83 0 2E-12
R132 98 1 250
I9 1 38 -1E-3
R133 5 58 1E9
D19 99 78 DD
X10 69 38 56 D560
X11 5 38 57 D560
X12 55 4 48 P450
M1 99 80 98 98 MSD
R146 44 15 0.03
R147 50 9 0.03
R148 52 24 0.03
R149 46 30 0.03
C30 4 6 1E-12
.MODEL DVN D KF=5E-16
.MODEL MSD PMOS KP=0.05 VTO=-2
.MODEL Q222 NPN IS=2E-13
.MODEL Q908 PNP IS=1E-13
.MODEL DD D
.MODEL DZ D BV=7.257 IBV=0.001 RS=5
.MODEL N912 NJF VTO=-3 BETA=3.2E-3 RS=12 RD=50
+ IS=1E-18 LAMBDA=3E-4 CGS=10E-12 CGD=0.5E-12
.MODEL C5V6 D IS=1E-15 RS=5 N=1 BV=5.6 IBV=1E-4
.MODEL C8V2 D IS=1E-15 RS=5 N=1 BV=8.2 IBV=1E-4
.MODEL Q907 PNP IS=1.1E-13 BF=150 BR=6 NF=1.2
+ RC=1 IKF=0.1 VAF=90 XTB=1.5 NE=1.8 ISE=1.5E-13
+ CJE=20E-12 VJE=0.8 MJE=1.2 CJC=15E-12 VJC=0.57
+ MJC=0.3 TF=0.5E-9 TR=35E-9
.ENDS MP230
.SUBCKT D560 10 20 30
M1 10 20 30 30 DMOS L=1U W=1U
CGS 20 30 43E-12
.MODEL DMOS NMOS LEVEL=3 VMAX=9E5 THETA=6E-3 ETA=2E-4
+ VTO=-2.5 KP=0.07 RS=2 RD=19
.ENDS
.SUBCKT P450 10 20 30
M1 10 20 30 30 DMOS L=1U W=1U
RDS 10 30 1E6
CGS 20 30 85E-12
CDG 10 20 20E-12
.MODEL DMOS PMOS LEVEL=3 VMAX=9E5 THETA=60E-3 ETA=2E-3
+ VTO=-2 KP=0.05 RS=3 RD=10
.ENDS
.SUBCKT irf540ns 1 2 3
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on Apr 24, 96
* Model format: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
* Default values used in MM:
* The voltage-dependent capacitances are
* not included. Other default values are:
*   RS=0 RD=0 LD=0 CBD=0 CBS=0 CGBO=0
.MODEL MM NMOS LEVEL=1 IS=1e-32
+VTO=3.55958 LAMBDA=0.000888191 KP=28.379
+CGSO=1.23576e-05 CGDO=1.77276e-08
RS 8 3 0.0251193
D1 3 1 MD
.MODEL MD D IS=1.13149e-09 RS=0.0078863 N=1.32265 BV=100
+IBV=0.00025 EG=1.17475 XTI=3.00167 TT=0
+CJO=7.95433e-10 VJ=0.5 M=0.374991 FC=0.5
RDS 3 1 4e+06
RD 9 1 0.00623556
RG 2 7 4.10175
D2 4 5 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=1.75616e-09 VJ=0.513551 M=0.614054 FC=1e-08
D3 0 5 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=3e-15 N=0.40002 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 3.86673e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=3e-15 N=0.40002
.ENDS
.SUBCKT irf9540n 1 2 3
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on Nov 20, 97
* MODEL FORMAT: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
* Default values used in MM:
* The voltage-dependent capacitances are
* not included. Other default values are:
*   RS=0 RD=0 LD=0 CBD=0 CBS=0 CGBO=0
.MODEL MM PMOS LEVEL=1 IS=1e-32
+VTO=-3.76841 LAMBDA=0 KP=7.07146
+CGSO=1.11762e-05 CGDO=1e-11
RS 8 3 0.0425484
D1 1 3 MD
.MODEL MD D IS=9.2473e-11 RS=0.00815502 N=1.22578 BV=100
+IBV=0.00025 EG=1.2 XTI=4 TT=6.92199e-07
+CJO=7.99077e-10 VJ=1.46806 M=0.554057 FC=0.499996
RDS 3 1 1e+06
RD 9 1 0.0462318
RG 2 7 7.07132
D2 5 4 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=2.43656e-09 VJ=1.23601 M=0.748171 FC=1e-08
D3 5 0 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=3e-15 N=0.4 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 3.41908e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 6 0 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=3e-15 N=0.4
.ENDS
* END MODEL MP230
***********
* REVISION 1 29-NOV-2005
* BEGIN MODEL MP240
* PINOUT ORDER +IN -IN +VB -VB GND CC1 CC2 IQ LSD HSD
*               41  42  1   38  2   6   4   5  7   8
*              +VS RS1 RS2 +ILIM -ILIM RS3 RS4 -VS
*               12  9   15   36    35   24  30  21
*
.SUBCKT MP240 41 42 1 38 2 6 4 5 7 8 12 9 15 36 35 24 30 21
X1 12 43 44 IRF640NS
X7 21 45 46 IRF9640
R77 47 1 39
C1 1 48 470E-12
X8 12 49 50 IRF640NS
X9 21 51 52 IRF9640
R82 53 49 10
R83 53 43 10
R84 54 51 10
R85 54 45 10
R86 6 55 100
R93 38 56 904
R94 38 57 278
Q12 4 47 1 Q907
D6 4 1 C8V2
E2 58 5 1 38 -30E-6
D8 59 0 DD
I1 0 59 1E-3
V16 59 60 0.7
E3 61 0 60 0 -571
R98 0 60 1E6
R99 0 61 1E6
E4 53 55 0 62 1.16E-3
E5 54 5 62 0 1.16E-3
V17 61 62 27
R100 0 62 1E6
D9 58 55 DZ
D10 63 64 C5V6
J2 63 65 66 N912
J3 4 67 68 N912
R101 69 66 51
R102 69 68 51
Q13 64 70 71 Q907
Q14 4 64 72 Q907
R103 71 1 200
R104 72 1 200
J4 4 63 4 N912
R105 63 64 1E5
D11 71 1 C8V2
V18 67 73 -4.0E-3
R106 64 70 70
C3 53 54 0.01E-6
R109 48 47 75
Q15 74 75 35 Q222
Q16 76 75 35 Q908
R110 75 36 100
Q17 76 52 77 Q908
R111 77 78 130
R112 77 79 5.1
Q18 74 78 79 Q222
R113 80 1 7000
Q20 80 8 81 Q222
R115 7 81 5600
D15 53 74 C5V6
D16 76 54 C5V6
R116 42 65 10
R117 41 82 10
C4 1 2 470E-12
C5 2 38 470E-12
E99 83 84 85 0 0.15
R118 85 86 1E6
R119 0 85 100
C25 86 85 1E-12
E100 86 0 1 0 1
R120 84 83 1E9
E101 84 87 88 0 0.15
R121 88 89 1E6
R122 0 88 100
C26 89 88 20E-12
E102 89 0 38 0 1
R123 87 84 1E9
E103 87 90 91 0 -0.15
R124 91 92 1E6
R125 0 91 100
C27 92 91 20E-12
E104 92 0 93 0 1
R126 90 87 1E9
E105 90 82 94 95 4
D17 94 0 DVN
I7 0 94 100E-6
D18 95 0 DVN
I8 0 95 100E-6
R127 82 90 1E9
E106 96 0 83 0 1
E107 97 0 65 0 1
R128 93 96 1E3
R129 93 97 1E3
R130 38 1 22E3
E108 73 83 62 0 40E-6
R131 83 73 1E9
C28 65 0 2E-12
C29 83 0 2E-12
R132 98 1 250
I9 1 38 -2.5E-3
R133 5 58 1E9
D19 99 78 DD
X10 5 38 57 D560
X11 69 38 56 D560
X12 55 4 48 P450
M1 99 80 98 98 MSD
R145 44 15 0.03
R146 50 9 0.03
R147 52 24 0.03
R148 46 30 0.03
C30 4 6 1E-12
.MODEL DVN D KF=5E-16
.MODEL DD D
.MODEL MSD PMOS KP=0.05 VTO=-2
.MODEL Q222 NPN IS=2E-13
.MODEL Q908 PNP IS=1E-13
.MODEL DZ D BV=7.870 IBV=0.001 RS=5
.MODEL N912 NJF VTO=-3 BETA=3.2E-3 RS=12 RD=50
+ IS=1E-18 LAMBDA=3E-4 CGS=10E-12 CGD=0.5E-12
.MODEL C5V6 D IS=1E-15 RS=5 N=1 BV=5.6 IBV=1E-4
.MODEL C8V2 D IS=1E-15 RS=5 N=1 BV=8.2 IBV=1E-4
.MODEL Q907 PNP IS=1.1E-13 BF=150 BR=6 NF=1.2
+ RC=1 IKF=0.1 VAF=90 XTB=1.5 NE=1.8 ISE=1.5E-13
+ CJE=20E-12 VJE=0.8 MJE=1.2 CJC=15E-12 VJC=0.57
+ MJC=0.3 TF=0.5E-9 TR=35E-9
.ENDS MP240
.SUBCKT D560 10 20 30
M1 10 20 30 30 DMOS L=1U W=1U
CGS 20 30 43E-12
.MODEL DMOS NMOS LEVEL=3 VMAX=9E5 THETA=6E-3 ETA=2E-4
+ VTO=-2.5 KP=0.07 RS=2 RD=19)
.ENDS
.SUBCKT P450 10 20 30
M1 10 20 30 30 DMOS L=1U W=1U
RDS 10 30 1E6
CGS 20 30 85E-12
CDG 10 20 20E-12
.MODEL DMOS PMOS LEVEL=3 VMAX=9E5 THETA=60E-3 ETA=2E-3
+ VTO=-2 KP=0.05 RS=3 RD=10)
.ENDS
.SUBCKT irf640ns 1 2 3
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on Feb 14, 02
* MODEL FORMAT: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
.MODEL MM NMOS LEVEL=1 IS=1e-32
+VTO=4.12428 LAMBDA=0.00426564 KP=7.74523
+CGSO=1.06e-05 CGDO=1e-10
RS 8 3 1e-05
D1 3 1 MD
.MODEL MD D IS=4.09854e-11 RS=0.00724292 N=1.17043 BV=200
+IBV=0.00025 EG=1.2 XTI=4 TT=0
+CJO=8e-10 VJ=1.41926 M=0.676432 FC=0.5
RDS 3 1 1e+06
RD 9 1 0.1
RG 2 7 1.35527
D2 4 5 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=1.5322e-09 VJ=1.34184 M=0.9 FC=1e-08
D3 0 5 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=3e-15 N=0.693912 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 2.19598e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=3e-15 N=0.693912
.ENDS
.SUBCKT irf9640 1 2 3
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on May 21, 96
* Model format: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
* Default values used in MM:
* The voltage-dependent capacitances are
* not included. Other default values are:
*   RS=0 RD=0 LD=0 CBD=0 CBS=0 CGBO=0
.MODEL MM PMOS LEVEL=1 IS=1e-32
+VTO=-3.8062 LAMBDA=0.0228396 KP=10.7224
+CGSO=1.09465e-05 CGDO=1e-11
RS 8 3 0.101556
D1 1 3 MD
.MODEL MD D IS=1e-17 RS=0.185714 N=1.5 BV=200
+IBV=0.00025 EG=1.2 XTI=4 TT=1e-07
+CJO=1.22255e-09 VJ=2.42988 M=0.605683 FC=0.493595
RDS 3 1 2e+06
RD 9 1 0.261579
RG 2 7 6.81119
D2 5 4 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=8.6947e-10 VJ=2.34088 M=0.9 FC=1e-08
D3 5 0 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=3e-15 N=0.402798 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 1.8148e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 6 0 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=3e-15 N=0.402798
.ENDS
* END MODEL MP240
***********
* REVISION 1 OCT-20-2006
* BEGIN MODEL MP38
* PINOUT ORDER +IN -IN +ILIM -ILIM OUT +VB -VB CC1 CC2 +VS -VS
*               29  30   24    23   15  1   26  6   4   12  18
.SUBCKT MP38 29 30 24 23 15 1 26 6 4 12 18
R77 31 1 20
C1 1 31 0.1E-6
X8 12 32 33 IRF640NS
X9 18 34 35 IRF9640
R82 36 32 51
R84 37 34 51
R86 6 38 100
R93 26 39 425
R94 26 40 157
Q12 4 31 1 Q907
D6 4 1 C8V2
E2 41 42 1 26 -30E-6
D8 43 0 DD
I1 0 43 1E-3
V16 43 44 0.7
E3 45 0 44 0 -571
R98 0 44 1E6
R99 0 45 1E6
E4 36 38 0 46 1.17E-3
E5 37 42 46 0 1.17E-3
V17 45 46 27
R100 0 46 1E6
D9 41 38 DZ
D10 47 48 C5V6
J2 47 49 50 N912
J3 4 51 52 N912
R101 53 50 30
R102 53 52 30
Q13 48 54 55 Q907C
Q14 4 48 56 Q907C
R103 55 1 100
R104 56 1 100
J4 4 47 4 N912
R105 47 48 1E5
D11 55 1 C8V2
V18 51 57 -1.5E-3
R106 48 54 160
C3 36 37 1E-9
Q15 58 59 23 Q222
Q16 37 59 23 Q908
R110 59 24 1
D15 36 58 C5V6
R116 30 49 51
R117 29 60 51
C4 1 61 470E-12
C5 61 26 470E-12
E99 62 63 64 0 0.15
R118 64 65 1E6
R119 0 64 100
C25 65 64 1E-12
E100 65 0 1 0 1
R120 63 62 1E9
E101 63 66 67 0 -0.15
R121 67 68 1E6
R122 0 67 100
C26 68 67 20E-12
E102 68 0 26 0 1
R123 66 63 1E9
E103 66 69 70 0 0.055
R124 70 71 1E6
R125 0 70 100
C27 71 70 20E-12
E104 71 0 72 0 1
R126 69 66 1E9
E105 69 60 73 74 4
D17 73 0 DVN
I7 0 73 100E-6
D18 74 0 DVN
I8 0 74 100E-6
R127 60 69 1E9
E106 75 0 62 0 1
E107 76 0 49 0 1
R128 72 75 1E3
R129 72 76 1E3
R130 26 1 100E3
E108 57 62 46 0 5E-6
R131 62 57 1E9
C28 49 0 2E-12
C29 62 0 2E-12
I9 1 26 -0.5E-3
R133 42 41 1E9
X10 53 26 39 D560
X11 42 26 40 D560
X12 38 4 31 P450
R141 0 61 1
R147 33 15 0.005
R148 35 15 0.12
.MODEL DVN D KF=5E-16
.MODEL MSD PMOS KP=0.05 VTO=-2
.MODEL Q222 NPN IS=2E-13
.MODEL Q908 PNP IS=1E-13
.MODEL DD D
.MODEL DZ D BV=7.833 IBV=0.001 RS=5
.MODEL N912 NJF VTO=-3 BETA=3.2E-3 RS=12 RD=50
+ IS=1E-18 LAMBDA=3E-4 CGS=10E-12 CGD=0.5E-12
.MODEL C5V6 D IS=1E-15 RS=5 N=1 BV=5.6 IBV=1E-4
.MODEL C8V2 D IS=1E-15 RS=5 N=1 BV=8.2 IBV=1E-4
.MODEL Q907 PNP IS=1.1E-13 BF=150 BR=6 NF=1.2
+ RC=1 IKF=0.1 VAF=90 XTB=1.5 NE=1.8 ISE=1.5E-13
+ CJE=20E-12 VJE=0.8 MJE=1.2 CJC=15E-12 VJC=0.57
+ MJC=0.3 TF=0.5E-9 TR=35E-9
.MODEL Q907C PNP IS=1.1E-13 BF=150 BR=6 NF=1.2
+ RC=1 IKF=0.1 VAF=500 XTB=1.5 NE=1.8 ISE=1.5E-13
+ CJE=20E-12 VJE=0.8 MJE=1.2 CJC=15E-12 VJC=0.57
+ MJC=0.3 TF=0.5E-9 TR=35E-9
.ENDS MP38
.SUBCKT D560 10 20 30
M1 10 20 30 30 DMOS L=1U W=1U
CGS 20 30 43E-12
.MODEL DMOS NMOS LEVEL=3 VMAX=9E5 THETA=6E-3 ETA=2E-4
+ VTO=-2.5 KP=0.07 RS=2 RD=19
.ENDS
.SUBCKT P450 10 20 30
M1 10 20 30 30 DMOS L=1U W=1U
RDS 10 30 1E6
CGS 20 30 85E-12
CDG 10 20 20E-12
.MODEL DMOS PMOS LEVEL=3 VMAX=9E5 THETA=60E-3 ETA=2E-3
+ VTO=-2 KP=0.05 RS=3 RD=10
.ENDS
.SUBCKT irf640ns 1 2 3
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on Feb 14, 02
* MODEL FORMAT: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
.MODEL MM NMOS LEVEL=1 IS=1e-32
+VTO=4.12428 LAMBDA=0.00426564 KP=7.74523
+CGSO=1.06e-05 CGDO=1e-10
RS 8 3 1e-05
D1 3 1 MD
.MODEL MD D IS=4.09854e-11 RS=0.00724292 N=1.17043 BV=200
+IBV=0.00025 EG=1.2 XTI=4 TT=0
+CJO=8e-10 VJ=1.41926 M=0.676432 FC=0.5
RDS 3 1 1e+06
RD 9 1 0.1
RG 2 7 1.35527
D2 4 5 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=1.5322e-09 VJ=1.34184 M=0.9 FC=1e-08
D3 0 5 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=3e-15 N=0.693912 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 2.19598e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=3e-15 N=0.693912
.ENDS
.SUBCKT irf9640 1 2 3
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on May 21, 96
* Model format: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
* Default values used in MM:
* The voltage-dependent capacitances are
* not included. Other default values are:
*   RS=0 RD=0 LD=0 CBD=0 CBS=0 CGBO=0
.MODEL MM PMOS LEVEL=1 IS=1e-32
+VTO=-3.8062 LAMBDA=0.0228396 KP=10.7224
+CGSO=1.09465e-05 CGDO=1e-11
RS 8 3 0.101556
D1 1 3 MD
.MODEL MD D IS=1e-17 RS=0.185714 N=1.5 BV=200
+IBV=0.00025 EG=1.2 XTI=4 TT=1e-07
+CJO=1.22255e-09 VJ=2.42988 M=0.605683 FC=0.493595
RDS 3 1 2e+06
RD 9 1 0.261579
RG 2 7 6.81119
D2 5 4 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=8.6947e-10 VJ=2.34088 M=0.9 FC=1e-08
D3 5 0 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=3e-15 N=0.402798 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 1.8148e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 6 0 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=3e-15 N=0.402798
.ENDS
* END MODEL MP38
************
* REVISION 1 OCT-20-2006
* BEGIN MODEL MP39
* PINOUT ORDER +IN -IN +ILIM -ILIM OUT +VB -VB CC1 CC2 +VS -VS
*               29  30   24    23   15  1   26  6   4   12  18
.SUBCKT MP39 29 30 24 23 15 1 26 6 4 12 18
R77 31 1 20
C1 1 31 0.1E-6
X8 12 32 33 IRF540NS
X9 18 34 35 IRF9540N
R82 36 32 51
R84 37 34 51
R86 6 38 100
R93 26 39 425
R94 26 40 157
Q12 4 31 1 Q907
D6 4 1 C8V2
E2 41 42 1 26 -5E-6
D8 43 0 DD
I1 0 43 1E-3
V16 43 44 0.7
E3 45 0 44 0 -571
R98 0 44 1E6
R99 0 45 1E6
E4 36 38 0 46 1.17E-3
E5 37 42 46 0 1.17E-3
V17 45 46 27
R100 0 46 1E6
D9 41 38 DZ
D10 47 48 C5V6
J2 47 49 50 N912
J3 4 51 52 N912
R101 53 50 30
R102 53 52 30
Q13 48 54 55 Q907C
Q14 4 48 56 Q907C
R103 55 1 100
R104 56 1 100
J4 4 47 4 N912
R105 47 48 1E5
D11 55 1 C8V2
V18 51 57 -1.5E-3
R106 48 54 160
C3 36 37 1E-9
Q15 58 59 23 Q222
Q16 37 59 23 Q908
R110 59 24 1
D15 36 58 C5V6
R116 30 49 51
R117 29 60 51
C4 1 61 470E-12
C5 61 26 470E-12
E99 62 63 64 0 0.15
R118 64 65 1E6
R119 0 64 100
C25 65 64 1E-12
E100 65 0 1 0 1
R120 63 62 1E9
E101 63 66 67 0 -0.15
R121 67 68 1E6
R122 0 67 100
C26 68 67 20E-12
E102 68 0 26 0 1
R123 66 63 1E9
E103 66 69 70 0 0.055
R124 70 71 1E6
R125 0 70 100
C27 71 70 20E-12
E104 71 0 72 0 1
R126 69 66 1E9
E105 69 60 73 74 4
D17 73 0 DVN
I7 0 73 100E-6
D18 74 0 DVN
I8 0 74 100E-6
R127 60 69 1E9
E106 75 0 62 0 1
E107 76 0 49 0 1
R128 72 75 1E3
R129 72 76 1E3
R130 26 1 100E3
E108 57 62 46 0 5E-6
R131 62 57 1E9
C28 49 0 2E-12
C29 62 0 2E-12
I9 1 26 -0.5E-3
R133 42 41 1E9
X10 53 26 39 D560
X11 42 26 40 D560
X12 38 4 31 P450
R141 0 61 1
R147 33 15 0.02
R148 35 15 0.05
.MODEL DVN D KF=5E-16
.MODEL MSD PMOS KP=0.05 VTO=-2
.MODEL Q222 NPN IS=2E-13
.MODEL Q908 PNP IS=1E-13
.MODEL DD D
.MODEL DZ D BV=7.228 IBV=0.001 RS=5
.MODEL N912 NJF VTO=-3 BETA=3.2E-3 RS=12 RD=50
+ IS=1E-18 LAMBDA=3E-4 CGS=10E-12 CGD=0.5E-12
.MODEL C5V6 D IS=1E-15 RS=5 N=1 BV=5.6 IBV=1E-4
.MODEL C8V2 D IS=1E-15 RS=5 N=1 BV=8.2 IBV=1E-4
.MODEL Q907 PNP IS=1.1E-13 BF=150 BR=6 NF=1.2
+ RC=1 IKF=0.1 VAF=90 XTB=1.5 NE=1.8 ISE=1.5E-13
+ CJE=20E-12 VJE=0.8 MJE=1.2 CJC=15E-12 VJC=0.57
+ MJC=0.3 TF=0.5E-9 TR=35E-9
.MODEL Q907C PNP IS=1.1E-13 BF=150 BR=6 NF=1.2
+ RC=1 IKF=0.1 VAF=500 XTB=1.5 NE=1.8 ISE=1.5E-13
+ CJE=20E-12 VJE=0.8 MJE=1.2 CJC=15E-12 VJC=0.57
+ MJC=0.3 TF=0.5E-9 TR=35E-9
.ENDS MP39
.SUBCKT D560 10 20 30
M1 10 20 30 30 DMOS L=1U W=1U
CGS 20 30 43E-12
.MODEL DMOS NMOS LEVEL=3 VMAX=9E5 THETA=6E-3 ETA=2E-4
+ VTO=-2.5 KP=0.07 RS=2 RD=19
.ENDS
.SUBCKT P450 10 20 30
M1 10 20 30 30 DMOS L=1U W=1U
RDS 10 30 1E6
CGS 20 30 85E-12
CDG 10 20 20E-12
.MODEL DMOS PMOS LEVEL=3 VMAX=9E5 THETA=60E-3 ETA=2E-3
+ VTO=-2 KP=0.05 RS=3 RD=10
.ENDS
.SUBCKT irf540ns 1 2 3
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on Apr 24, 96
* Model format: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
* Default values used in MM:
* The voltage-dependent capacitances are
* not included. Other default values are:
*   RS=0 RD=0 LD=0 CBD=0 CBS=0 CGBO=0
.MODEL MM NMOS LEVEL=1 IS=1e-32
+VTO=3.55958 LAMBDA=0.000888191 KP=28.379
+CGSO=1.23576e-05 CGDO=1.77276e-08
RS 8 3 0.0251193
D1 3 1 MD
.MODEL MD D IS=1.13149e-09 RS=0.0078863 N=1.32265 BV=100
+IBV=0.00025 EG=1.17475 XTI=3.00167 TT=0
+CJO=7.95433e-10 VJ=0.5 M=0.374991 FC=0.5
RDS 3 1 4e+06
RD 9 1 0.00623556
RG 2 7 4.10175
D2 4 5 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=1.75616e-09 VJ=0.513551 M=0.614054 FC=1e-08
D3 0 5 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=3e-15 N=0.40002 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 3.86673e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=3e-15 N=0.40002
.ENDS
.SUBCKT irf9540n 1 2 3
**************************************
*      Model Generated by MODPEX     *
*Copyright(c) Symmetry Design Systems*
*         All Rights Reserved        *
*    UNPUBLISHED LICENSED SOFTWARE   *
*   Contains Proprietary Information *
*      Which is The Property of      *
*     SYMMETRY OR ITS LICENSORS      *
*Commercial Use or Resale Restricted *
*   by Symmetry License Agreement    *
**************************************
* Model generated on Nov 20, 97
* MODEL FORMAT: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
* Default values used in MM:
* The voltage-dependent capacitances are
* not included. Other default values are:
*   RS=0 RD=0 LD=0 CBD=0 CBS=0 CGBO=0
.MODEL MM PMOS LEVEL=1 IS=1e-32
+VTO=-3.76841 LAMBDA=0 KP=7.07146
+CGSO=1.11762e-05 CGDO=1e-11
RS 8 3 0.0425484
D1 1 3 MD
.MODEL MD D IS=9.2473e-11 RS=0.00815502 N=1.22578 BV=100
+IBV=-0.00025 EG=1.2 XTI=4 TT=6.92199e-07
+CJO=7.99077e-10 VJ=1.46806 M=0.554057 FC=0.499996
RDS 3 1 1e+06
RD 9 1 0.0462318
RG 2 7 7.07132
D2 5 4 MD1
* Default values used in MD1:
*   RS=0 EG=1.11 XTI=3.0 TT=0
*   BV=infinite IBV=1mA
.MODEL MD1 D IS=1e-32 N=50
+CJO=2.43656e-09 VJ=1.23601 M=0.748171 FC=1e-08
D3 5 0 MD2
* Default values used in MD2:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   BV=infinite IBV=1mA
.MODEL MD2 D IS=3e-15 N=0.4 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 3.41908e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 6 0 MD3
* Default values used in MD3:
*   EG=1.11 XTI=3.0 TT=0 CJO=0
*   RS=0 BV=infinite IBV=1mA
.MODEL MD3 D IS=3e-15 N=0.4
.ENDS
* END MODEL MP39
**********
*REVISION 3 26-NOV-2004
*REVISED GAIN AND PHASE TO MATCH NEW DATA SHEET
*MADE ILIMIT SYMMETRIC, ADJUSTED IQ
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA01
* BEGIN OPAMP MACROMODEL PA01
* PINOUT ORDER +IN -IN RCL+ RCLC RCL- OUT +V -V
*                1   2  29   31   30   3   4  5
.SUBCKT PA01 1 2 29 31 30 3 4 5
* POSITIVE CURRENT LIMIT RESISTOR GOES FROM RCL+ TO RCLC
* NEGATIVE CURRENT LIMIT RESISTOR GOES FROM RCL- TO RCLC
* NOTE THAT CURRENT LIMIT RESISTORS DO NOT CONNECT TO THE OUTPUT
* LIKE THEY DO IN THE PHYSICAL PART
Q1 10 1 8 QI1
Q2 11 2 9 QI2
R3 12 8 2.68E+03
R4 12 9 2.68E+03
I2 12 5 3.10E-05
C1 12 5 1.43E-12
R5 12 5 2.50E+08
R1 4 10 3.98E+03
R2 4 11 3.98E+03
C2 10 11 5E-12
I1 4 5 9.7E-03
G1 6 0 11 10 2.51E-04
G2 6 0 12 0 1.41E-09
R6 6 0 1.00E+05
D1 6 0 DD
D2 0 6 DD
C3 6 7 1E-11
G3 0 7 0 6 4.50E+00
R7 7 0 1E3
D3 7 16 DD
V1 18 16 5.70E+00
D4 17 7 DD
V2 17 19 5.70E+00
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 0 2.78E-10
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 1.08E-01
R13 22 24 1.08E-01
D5 23 25 DL
D6 26 24 DL
R9 27 29 550
R10 28 30 550
I3 18 23 9.93E-03
I4 24 19 9.93E-03
R15 31 3 6.67E-01
DC1 3 4 DO
DC2 5 3 DO
.MODEL DO D(CJO=10PF IS=5.77E-14 RS=5.19E-02)
RS1 29 31 1E6
RS2 30 31 1E6
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL QI1 NPN (BF=2.29E+03 IS=8E-16)
.MODEL QI2 NPN (BF=1.63E+03 IS=9.54E-16)
.MODEL QOP PNP (BF=5.82E+02 IS=1E-14)
.MODEL QON NPN (BF=5.82E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-12)
.MODEL QLP PNP (BF=100 IS=1E-12)
* END OF OPAMP MACROMODEL
.ENDS
***********
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA01
* BEGIN OPAMP MACROMODEL PA02
* PINOUT ORDER +IN -IN RCL+ RCLC RCL- OUT +V -V
*                1   2  29   31   30   3   4  5
.SUBCKT PA02 1 2 29 31 30 3 4 5
* POSITIVE CURRENT LIMIT RESISTOR GOES FROM RCL+ TO RCLC
* NEGATIVE CURRENT LIMIT RESISTOR GOES FROM RCL- TO RCLC
* NOTE THAT CURRENT LIMIT RESISTORS DO NOT CONNECT TO THE SUPPLIES
* LIKE THEY DO IN THE PHYSICAL PART
J1 10 1 8 JI1
J2 11 2 9 JI2
R3 12 8 1.52E+03
R4 12 9 1.52E+03
I2 12 5 1.00E-04
C1 12 5 5.56E-13
R5 12 5 4.00E+07
R1 4 10 1.77E+03
R2 4 11 1.77E+03
C2 10 11 9.00E-12
I1 4 5 1.74E-02
G1 6 15 11 10 5.65E-04
G2 6 15 12 15 1.79E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 5.00E-12
G3 15 7 15 6 2.50E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 1.20E+00
D4 17 7 DD
V2 17 19 1.20E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 3.12E-11
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 1.19E-01
R13 22 24 1.19E-01
D5 23 25 DL
D6 26 24 DL
R9 27 29 1E3
R10 28 30 100
I3 18 23 9.47E-03
I4 24 19 9.47E-03
R15 31 3 4.18E-01
DC1 3 4 DO
DC2 5 3 DO
.MODEL DO D(CJO=10PF IS=5.25E-14 RS=5.71E-02)
RS1 29 31 1E6
RS2 30 31 1E6
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL JI1 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1)
.MODEL JI2 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1.0050)
.MODEL QOP PNP (BF=5.54E+02 IS=1E-14)
.MODEL QON NPN (BF=5.54E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
**********
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA09
* BEGIN OPAMP MACROMODEL PA03
* PINOUT ORDER +IN -IN OUT +V -V COMP COMP
*                1   2  3   4  5   6    7
.SUBCKT PA03 1 2 3 4 5 6 7
J1 10 1 8 JI1
J2 11 2 9 JI2
R3 12 8 5.08E+02
R4 12 9 5.08E+02
I2 12 5 9.00E-04
C1 12 5 7.00E-12
R5 12 5 1.79E+06
R1 4 10 7.58E+02
R2 4 11 7.58E+02
C2 10 11 1.75E-10
I1 4 5 9.95E-02
G1 6 15 11 10 1.32E-03
G2 6 15 12 15 7.42E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 100E-12
G3 15 7 15 6 2.40E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 3.20E+00
D4 17 7 DD
V2 17 19 3.20E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 9.19E-10
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 1.75E-02
RCLP 29 31 1.75E-02
RCLN 30 31 1.75E-02
R13 22 24 1.75E-02
D5 23 25 DL
D6 26 24 DL
R9 27 29 1E3
R10 28 30 1E3
I3 18 23 2.47E-02
I4 24 19 2.47E-02
R15 31 3 1.17E-01
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=3.57E-13 RS=8.40E-03)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL JI1 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1)
.MODEL JI2 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1.0005)
.MODEL QOP PNP (BF=1.45E+03 IS=1E-14)
.MODEL QON NPN (BF=1.45E+03 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
**********
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*ADDED BUFFER STAGE BETWEEN INPUT & OUTPUT
*SYM=PA04
* BEGIN OPAMP MACROMODEL PA04
* PINOUT ORDER  +IN -IN OUT ILIM-10 ILIM-11 +VB -VB COMP COMP +VS -VS
*                 1   2  3    33      31     4    5   6    7   36  37
.SUBCKT PA04 1 2 3 33 31 4 5 6 7 36 37
M1 10 1 8 8 MI1
M2 11 2 9 9 MI2
R3 12 8 5.00E+01
R4 12 9 5.00E+01
I2 12 5 6.65E-03
C1 12 5 7.92E-11
R5 12 5 3.01E+06
R1 4 10 8.38E+01
R2 4 11 8.38E+01
C2 10 11 1.90E-10
I1 4 5 2.18E-02
G1 6 15 11 10 1.19E-02
G2 6 15 12 15 3.77E-08
R6 6 15 6.21E+04
D1 6 34 DD
D7 34 15 DD
D2 35 6 DD
D8 15 35 DD
C3 6 7 33.0E-12
G3 15 7 15 6 1.35E-01
R7 7 15 1E3
D3 7 16 DD
V1 18 16 5.95E+00
D4 17 7 DD
V2 17 19 5.95E+00
RE1 15 0 0.001
E2 38 0 4 0 1
E3 39 0 5 0 1
R8 7 20 50
C4 20 15 1.42E-10
Q3 37 20 21 QOP
Q4 36 20 22 QON
Q5 36 21 29 QON
Q6 37 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 31 1E3
R10 28 31 1E3
E4 41 36 38 36 0.65
E5 42 37 39 37 0.65
E6 18 0 41 0 1
E7 19 0 42 0 1
RY1 38 0 10E6
RY2 39 0 10E6
RY3 39 0 10E6
RY4 41 0 10E6
I3 36 21 1.99E-02
I4 22 37 1.99E-02
R15 29 3 2.25E-01
DC1 29 36 DO
DC2 37 29 DO
I5 37 36 1.97E-02
.MODEL DO D(CJO=10PF IS=2.31E-13 RS=1.30E-02)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MI1 NMOS (KP=2.96E-02 IS=3E-16 VTO=1)
.MODEL MI2 NMOS (KP=2.96E-02 IS=3E-16 VTO=0.9950)
.MODEL QOP PNP (BF=1.16E+03 IS=1E-14)
.MODEL QON NPN (BF=1.16E+03 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*ADDED BURRER BETWEEN INPUT AND OUTPUT
*SYM=PA04
* BEGIN OPAMP MACROMODEL PA05
* PINOUT ORDER  +IN -IN OUT ILIM-10 ILIM-11 +VB -VB
* PINOUT ORDER CONTINUED  COMP COMP +VS -VS
.SUBCKT PA05 1 2 3 33 31 4 5 6 7 36 37
M1 10 1 8 8 MI1
M2 11 2 9 9 MI2
R3 12 8 5.40E+01
R4 12 9 5.40E+01
I2 12 5 8.99E-03
C1 12 5 1.76E-12
R5 12 5 2.76E+06
R1 4 10 1.26E+02
R2 4 11 1.26E+02
C2 10 11 2.10E-10
I1 4 5 3.69E-02
G1 6 15 11 10 7.91E-03
G2 6 15 12 15 7.91E-08
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 5.00E-12
G3 15 7 15 6 1.59E-01
R7 7 15 1E3
D3 7 16 DD
V1 18 16 6.70E+00
D4 17 7 DD
V2 17 19 6.70E+00
RE1 15 0 0.001
E2 38 0 4 0 1
E3 39 0 5 0 1
R8 7 20 50
C4 20 15 3.79E-10
Q3 37 20 21 QOP
Q4 36 20 22 QON
Q5 36 21 29 QON
Q6 37 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 31 1E3
R10 28 31 1E3
E4 41 36 38 36 1
E5 42 37 39 37 1
E6 18 0 41 0 1
E7 19 0 42 0 1
RY1 38 0 10E6
RY2 39 0 10E6
RY3 41 0 10E6
RY4 42 0 10E6
I3 36 21 7.15E-03
I4 22 37 7.15E-03
R15 29 3 1.58E-01
DC1 29 36 DO
DC2 37 29 DO
I5 36 37 2.25E-02
.MODEL DO D(CJO=10PF IS=3.99E-13 RS=7.52E-03)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MI1 NMOS (KP=1.38E-02 IS=3E-16 VTO=1)
.MODEL MI2 NMOS (KP=1.38E-02 IS=3E-16 VTO=0.9950)
.MODEL QOP PNP (BF=5.58E+03 IS=1E-14)
.MODEL QON NPN (BF=5.58E+03 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
**************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA01
* BEGIN OPAMP MACROMODEL PA07
* PINOUT ORDER +IN -IN RCL+ RCLC RCL- OUT +V -V
*                1   2  29   31   30   3   4  5
.SUBCKT PA07 1 2 29 31 30 3 4 5
* POSITIVE CURRENT LIMIT RESISTOR GOES FROM RCL+ TO RCLC
* NEGATIVE CURRENT LIMIT RESISTOR GOES FROM RCL- TO RCLC
* NOTE THAT CURRENT LIMIT RESISTORS DO NOT CONNECT TO THE OUTPUT
* LIKE THEY DO IN THE PHYSICAL PART
J1 10 1 8 JI1
J2 11 2 9 JI2
R3 12 8 1.57E+04
R4 12 9 1.57E+04
I2 12 5 2.50E-05
C1 12 5 2.08E-13
R5 12 5 4.00E+07
R1 4 10 1.59E+04
R2 4 11 1.59E+04
C2 10 11 2.50E-12
I1 4 5 8.04E-03
G1 6 15 11 10 6.28E-05
G2 6 15 12 15 6.28E-11
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 5.00E-12
G3 15 7 15 6 1.59E+01
R7 7 15 1E3
D3 7 16 DD
V1 18 16 3.70E+00
D4 17 7 DD
V2 17 19 3.70E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 9.17E-11
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 1.08E-01
R13 22 24 1.08E-01
D5 23 25 DL
D6 26 24 DL
R9 27 29 1E3
R10 28 30 100
I3 18 23 9.93E-03
I4 24 19 9.93E-03
R15 31 3 3.25E-01
DC1 3 4 DO
DC2 5 3 DO
.MODEL DO D(CJO=10PF IS=5.77E-14 RS=5.19E-02)
RS1 29 31 1E6
RS2 30 31 1E6
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL JI1 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1)
.MODEL JI2 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1.0005)
.MODEL QOP PNP (BF=5.82E+02 IS=1E-14)
.MODEL QON NPN (BF=5.82E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
******************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA01
* BEGIN OPAMP MACROMODEL PA08
* PINOUT ORDER +IN -IN RCL+ RCLC RCL- OUT +V -V
*                1   2  29   31   30   3   4  5
.SUBCKT PA08 1 2 29 31 30 3 4 5
* POSITIVE CURRENT LIMIT RESISTOR GOES FROM RCL+ TO RCLC
* NEGATIVE CURRENT LIMIT RESISTOR GOES FROM RCL- TO RCLC
* NOTE THAT CURRENT LIMIT RESISTORS DO NOT CONNECT TO THE OUTPUT
* LIKE THEY DO IN THE PHYSICAL PART
J1 10 1 8 JI1
J2 11 2 9 JI2
R3 12 8 2.40E+03
R4 12 9 2.40E+03
I2 12 5 1.50E-04
C1 12 5 3.57E-13
R5 12 5 2.00E+08
R1 4 10 2.65E+03
R2 4 11 2.65E+03
C2 10 11 4.29E-12
I1 4 5 4.08E-03
G1 6 15 11 10 3.77E-04
G2 6 15 12 15 1.19E-10
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 5.00E-12
G3 15 7 15 6 1.49E+01
R7 7 15 1E3
D3 7 16 DD
V1 18 16 3.70E+00
D4 17 7 DD
V2 17 19 3.70E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 2.22E-11
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 3.40E+00
R13 22 24 3.40E+00
D5 23 25 DL
D6 26 24 DL
R9 27 29 1E3
R10 28 30 100
I3 18 23 1.77E-03
I4 24 19 1.77E-03
R15 31 3 3.57E+01
RS1 29 31 1E6
RS2 30 31 1E6
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL JI1 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1)
.MODEL JI2 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1.0005)
.MODEL QOP PNP (BF=1.04E+02 IS=1E-14)
.MODEL QON NPN (BF=1.04E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
**********************
* REVISION 3 1/13/2003
* SYM=PA09
* MAJOR CHANGE TO REFLECT DATA SHEET CHANGES OF
* JANUARY 2003.  THIS MODEL DOES NOT FOLLOW
* LARGE SIGNAL PERFORMANCE IN THE FOLLOWING AREAS:
*   QUIESCENT DOES NOT INCREASE WITH HIGH DV/DT SIGNALS.
*   PHASE MARGIN DOES NOT MOVE WITH SUPPLIES, SWING
*   TO THE RAIL, OR LOADING.
*   DOES NOT SHOW OVERLOAD RECOVERY TIME.
* WHILE THIS MODEL ACCURATELY REPRESENTS SMALL SIGNAL
* PARAMETERS, SLEW RATE AND OUTPUT IMPEDANCE, IT IS
* RECOMMENDED THAT THE HARDWARE BE TESTED WITH THE 
* TECHNIQUE PRESENTED IN AP NOTE 19, FIGURES 40 AND 41.
* EXPAND THIS TEST TO LARGE SIGNAL LEVELS TO REVEAL
* POSSIBLE PROBLEMS THIS MODEL WILL NOT SHOW.
* BEGIN OPAMP MACROMODEL PA09
* PINOUT ORDER +IN -IN OUT +V -V COMP COMP
*               1   2   3   4  5   6    7
.SUBCKT PA09 1 2 3 4 5 6 7
J1 10 1 8 JI1
J2 11 2 9 JI2
R3 12 8 350
R4 12 9 350
C8 8 9 10E-12
I2 12 5 4.20E-03
C1 12 5 4.57E-14
R5 12 5 2.00E+06
R1 4 10 66.3
R2 4 11 66.3
C2 10 11 1.33E-10
I1 4 5 6.59E-02
G1 6 15 11 10 3.00E-02
G2 6 15 12 15 9.51E-08
R6 6 15 1.10E+05
D1 6 34 DD
D7 34 15 DD
D2 35 6 DD
D8 15 35 DD
C3 6 7 2.50E-13
G3 15 7 15 6 14.35E-02
R7 7 15 1E3
D3 7 16 DD
V1 18 16 6.70E+00
D4 17 7 DD
V2 17 19 6.70E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 50 120.5
C4 50 15 3.65E-11
E50 51 0 50 0 1
E60 61 0 50 0 1
D50 7 61 DD
D51 61 7 DD
R58 51 20 50
C54 20 15 262E-12
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 7.44E-02
RCLP 29 31 7.44E-02
RCLN 30 31 7.44E-02
R13 22 24 7.44E-02
D5 23 25 DL
D6 26 24 DL
R9 27 29 1E3
R10 28 30 1E3
I3 18 23 1.86E-03
I4 24 19 1.86E-03
R15 31 3 5.00E-01
DC1 31 4 DO
DC2 5 31 DO
.MODEL DO D(CJO=10PF IS=8.40E-14 RS=3.57E-02)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL JI1 NJF (BETA=6.35E-02 IS=3E-16 VTO=-1)
.MODEL JI2 NJF (BETA=6.35E-02 IS=3E-16 VTO=-1.0030)
.MODEL QOP PNP (BF=4.52E+03 IS=1E-14)
.MODEL QON NPN (BF=4.52E+03 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
*************
*REVISION 3 25-NOV-2004
*CHANGED GAIN AND PHASE TO MATCH BENCH DATA
*ADJUSTED IQ AND VDROP TO MATCH DATA SHEET
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY
*SYM=PA10
* BEGIN OPAMP MACROMODEL PA10
* PINOUT ORDER +IN -IN OUT +V -V CL+ CL- FO
*                1   2  3   4  5  35 36  37
.SUBCKT PA10 1 2 3 4 5 35 36 37
Q1 10 1 8 QI1
Q2 11 2 9 QI2
R3 12 8 2.68E+03
R4 12 9 2.68E+03
I2 12 5 3.10E-05
C1 12 5 1.43E-12
R5 12 5 2.50E+08
R1 4 10 3.98E+03
R2 4 11 3.98E+03
C2 10 11 5E-12
I1 4 5 1.5E-03
G1 6 0 11 10 2.51E-04
G2 6 0 12 0 1.41E-09
R6 6 0 1.00E+05
D1 6 0 DD
D2 0 6 DD
C3 6 7 1.00E-11
G3 0 7 0 6 4.5E+00
R7 7 0 1E3
D3 7 16 DD
V1 18 16 3E+00
D4 17 7 DD
V2 17 19 4.50E+00
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 0 278E-12
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 3 QLN
Q8 26 28 3 QLP
R11 21 23 3.97E-02
RF1 27 37 20E3
RF2 28 37 20E3
R13 22 24 3.97E-02
D5 23 25 DL
D6 26 24 DL
R9 27 35 280
R10 28 36 280
I3 18 23 1.64E-02
I4 24 19 1.64E-02
RO1 29 35 0.402
RO2 30 36 0.402
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL QI1 NPN (BF=2.22E+03 IS=8E-16)
.MODEL QI2 NPN (BF=1.33E+03 IS=8.62E-16)
.MODEL QOP PNP (BF=3.20E+02 IS=1E-14)
.MODEL QON NPN (BF=3.20E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=4E-13)
.MODEL QLP PNP (BF=100 IS=4E-13)
* END OF OPAMP MACROMODEL
.ENDS
*****************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA10
* BEGIN OPAMP MACROMODEL PA12
* PINOUT ORDER +IN -IN OUT +V -V CL+ CL- FO
*                1   2  3   4  5  35 36  37
.SUBCKT PA12 1 2 3 4 5 35 36 37
Q1 10 1 8 QI1
Q2 11 2 9 QI2
R3 12 8 2.68E+03
R4 12 9 2.68E+03
I2 12 5 4.00E-05
C1 12 5 1.43E-12
R5 12 5 2.50E+07
R1 4 10 3.98E+03
R2 4 11 3.98E+03
C2 10 34 15E-12
RZ 34 11 40
I1 4 5 8.56E-03
G1 6 15 11 10 2.51E-04
G2 6 15 12 15 1.41E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 1.00E-11
G3 15 7 15 6 7.08E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 2.70E+00
D4 17 7 DD
V2 17 19 4.50E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 1E-12
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 3 QLNA
Q8 26 28 3 QLPA
R11 21 23 3.97E-02
RF1 27 37 20E3
RF2 28 37 20E3
R13 22 24 3.97E-02
D5 23 25 DL
D6 26 24 DL
R9 27 35 280
R10 28 36 280
I3 18 23 1.64E-02
I4 24 19 1.64E-02
RO1 29 35 0.134
RO2 30 36 0.134
RFF1 37 35 10E6
RFF2 37 36 10E6
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL QI1 NPN (BF=2.22E+03 IS=8E-16)
.MODEL QI2 NPN (BF=1.33E+03 IS=8.62E-16)
.MODEL QOP PNP (BF=9.60E+02 IS=1E-14)
.MODEL QON NPN (BF=9.60E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
.MODEL QLNA NPN (BF=100 IS=4E-13)
.MODEL QLPA PNP (BF=100 IS=4E-13)
* END OF OPAMP MACROMODEL
.ENDS
*******************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA10
* BEGIN OPAMP MACROMODEL PA13
* PINOUT ORDER +IN -IN OUT +V -V CL+ CL- FO
*                1   2  3   4  5  35 36  37
.SUBCKT PA13 1 2 3 4 5 35 36 37
Q1 10 1 8 QI1
Q2 11 2 9 QI2
R3 12 8 2.68E+03
R4 12 9 2.68E+03
I2 12 5 4.00E-05
C1 12 5 1.43E-12
R5 12 5 2.50E+07
R1 4 10 3.98E+03
R2 4 11 3.98E+03
C2 10 34 15E-12
RZ 34 11 40
I1 4 5 8.56E-03
G1 6 15 11 10 2.51E-04
G2 6 15 12 15 1.41E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 1.00E-11
G3 15 7 15 6 7.08E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 2.70E+00
D4 17 7 DD
V2 17 19 4.50E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 1E-12
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 3 QLNA
Q8 26 28 3 QLPA
R11 21 23 3.97E-02
RF1 27 37 20E3
RF2 28 37 20E3
R13 22 24 3.97E-02
D5 23 25 DL
D6 26 24 DL
R9 27 35 280
R10 28 36 280
I3 18 23 1.64E-02
I4 24 19 1.64E-02
RO1 29 35 0.134
RO2 30 36 0.134
RFF1 37 35 10E6
RFF2 37 36 10E6
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL QI1 NPN (BF=2.22E+03 IS=8E-16)
.MODEL QI2 NPN (BF=1.33E+03 IS=8.62E-16)
.MODEL QOP PNP (BF=9.60E+02 IS=1E-14)
.MODEL QON NPN (BF=9.60E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
.MODEL QLNA NPN (BF=100 IS=4E-13)
.MODEL QLPA PNP (BF=100 IS=4E-13)
* END OF OPAMP MACROMODEL
.ENDS
************
*REVISION 2 18-MAR-2002 RENAMED FROM PA40
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA09
* BEGIN OPAMP MACROMODEL PA140
* PINOUT ORDER +IN -IN OUT +V -V COMP COMP
*                1   2  3   4  5   6    7
.SUBCKT PA140 1 2 3 4 5 6 7
M1 10 1 8 8 MI1
M2 11 2 9 9 MI2
R3 12 8 2.95E+03
R4 12 9 2.95E+03
I2 12 5 2.90E-04
C1 12 5 7.78E-13
R5 12 5 1.38E+08
R1 4 10 3.20E+03
R2 4 11 3.20E+03
C2 10 11 1.66E-11
I1 4 5 -8.81E-05
G1 6 15 11 10 3.13E-04
G2 6 15 12 15 5.56E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 5.00E-12
G3 15 7 15 6 5.69E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 3.20E+00
D4 17 7 DD
V2 17 19 6.70E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 9.35E-11
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
M3 25 27 3 3 MLN
M4 26 28 3 3 MLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 1.20E-03
I4 22 19 1.20E-03
R15 29 3 7.50E+01
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=8.40E-16 RS=3.57E+00)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MI1 NMOS (KP=4.00E-03 IS=3E-16 VTO=1)
.MODEL MI2 NMOS (KP=4.00E-03 IS=3E-16 VTO=0.9850)
.MODEL MLN NMOS (KP=5.00E-03 IS=3E-16 VTO=2.5)
.MODEL MLP PMOS (KP=5.00E-03 IS=3E-16 VTO=-2.5)
.MODEL QOP PNP (BF=7.01E+01 IS=1E-14)
.MODEL QON NPN (BF=7.01E+01 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
************
*REVISION 2 18-MAR-2002 COPIED FROM PA41
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA85
* BEGIN OPAMP MACROMODEL PA141
* PINOUT ORDER +IN -IN CL OUT +V -V COMP COMP
*                1   2  3  33  4  5   6    7
.SUBCKT PA141 1 2 3 33 4 5 6 7
M1 10 1 8 8 MI1
M2 11 2 9 9 MI2
R3 12 8 2.95E+03
R4 12 9 2.95E+03
I2 12 5 2.90E-04
C1 12 5 7.78E-13
R5 12 5 1.38E+08
R1 4 10 3.20E+03
R2 4 11 3.20E+03
C2 10 11 1.66E-11
I1 4 5 -8.81E-05
G1 6 15 11 10 3.13E-04
G2 6 15 12 15 5.56E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 5.00E-12
G3 15 7 15 6 5.69E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 3.20E+00
D4 17 7 DD
V2 17 19 6.70E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 9.35E-11
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
M3 25 27 33 33 MLN
M4 26 28 33 33 MLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 1.20E-03
I4 22 19 1.20E-03
R15 29 3 7.50E+01
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=8.40E-16 RS=3.57E+00)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MI1 NMOS (KP=4.00E-03 IS=3E-16 VTO=1)
.MODEL MI2 NMOS (KP=4.00E-03 IS=3E-16 VTO=0.9850)
.MODEL MLN NMOS (KP=5.00E-03 IS=3E-16 VTO=2.5)
.MODEL MLP PMOS (KP=5.00E-03 IS=3E-16 VTO=-2.5)
.MODEL QOP PNP (BF=7.01E+01 IS=1E-14)
.MODEL QON NPN (BF=7.01E+01 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
*************
*REVISION 2 18-MAR-2002 COPIED FROM PA42
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA85
* BEGIN OPAMP MACROMODEL PA142
* PINOUT ORDER +IN -IN CL OUT +V -V COMP COMP
*                1   2  3  33  4  5   6    7
.SUBCKT PA142 1 2 3 33 4 5 6 7
M1 10 1 8 8 MI1
M2 11 2 9 9 MI2
R3 12 8 2.95E+03
R4 12 9 2.95E+03
I2 12 5 2.90E-04
C1 12 5 7.78E-13
R5 12 5 1.38E+08
R1 4 10 3.20E+03
R2 4 11 3.20E+03
C2 10 11 1.66E-11
I1 4 5 -8.81E-05
G1 6 15 11 10 3.13E-04
G2 6 15 12 15 5.56E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 5.00E-12
G3 15 7 15 6 5.69E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 3.20E+00
D4 17 7 DD
V2 17 19 6.70E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 9.35E-11
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
M3 25 27 33 33 MLN
M4 26 28 33 33 MLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 1.20E-03
I4 22 19 1.20E-03
R15 29 3 7.50E+01
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=8.40E-16 RS=3.57E+00)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MI1 NMOS (KP=4.00E-03 IS=3E-16 VTO=1)
.MODEL MI2 NMOS (KP=4.00E-03 IS=3E-16 VTO=0.9850)
.MODEL MLN NMOS (KP=5.00E-03 IS=3E-16 VTO=2.5)
.MODEL MLP PMOS (KP=5.00E-03 IS=3E-16 VTO=-2.5)
.MODEL QOP PNP (BF=7.01E+01 IS=1E-14)
.MODEL QON NPN (BF=7.01E+01 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
*************
*REVISION 2 18-MAR-2002 COPIED FROM PA44
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA85
* BEGIN OPAMP MACROMODEL PA144
* PINOUT ORDER +IN -IN CL OUT +V -V COMP COMP
*                1   2  3  33  4  5   6    7
.SUBCKT PA144 1 2 3 33 4 5 6 7
M1 10 1 8 8 MI1
M2 11 2 9 9 MI2
R3 12 8 2.95E+03
R4 12 9 2.95E+03
I2 12 5 2.90E-04
C1 12 5 7.78E-13
R5 12 5 1.38E+08
R1 4 10 3.20E+03
R2 4 11 3.20E+03
C2 10 11 1.66E-11
I1 4 5 -8.81E-05
G1 6 15 11 10 3.13E-04
G2 6 15 12 15 5.56E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 5.00E-12
G3 15 7 15 6 5.69E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 3.20E+00
D4 17 7 DD
V2 17 19 6.70E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 9.35E-11
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
M3 25 27 33 33 MLN
M4 26 28 33 33 MLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 1.20E-03
I4 22 19 1.20E-03
R15 29 3 7.50E+01
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=8.40E-16 RS=3.57E+00)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MI1 NMOS (KP=4.00E-03 IS=3E-16 VTO=1)
.MODEL MI2 NMOS (KP=4.00E-03 IS=3E-16 VTO=0.9850)
.MODEL MLN NMOS (KP=5.00E-03 IS=3E-16 VTO=2.5)
.MODEL MLP PMOS (KP=5.00E-03 IS=3E-16 VTO=-2.5)
.MODEL QOP PNP (BF=7.01E+01 IS=1E-14)
.MODEL QON NPN (BF=7.01E+01 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
*******************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA85
* BEGIN OPAMP MACROMODEL PA15
* PINOUT ORDER +IN -IN CL OUT +V -V COMP COMP
*                1   2  3  33  4  5   6    7
.SUBCKT PA15 1 2 3 33 4 5 6 7
M1 10 1 8 8 MI1
M2 11 2 9 9 MI2
R3 12 8 3.07E+03
R4 12 9 3.07E+03
I2 12 5 8.00E-05
C1 12 5 2.86E-12
R5 12 5 6.88E+07
R1 4 10 3.32E+03
R2 4 11 3.32E+03
C2 10 11 3.00E-12
I1 4 5 -3.99E-04
G1 6 15 11 10 5.21E-04
G2 6 15 12 15 3.79E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 5.00E-12
G3 15 7 15 6 1.87E+01
R7 7 15 1E3
D3 7 16 DD
V1 18 16 4.50E+00
D4 17 7 DD
V2 17 19 4.50E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 2.32E-09
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 4.32E-03
I4 22 19 1.72E-03
R15 29 3 5
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=3.15E-15 RS=9.52E-01)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MI1 NMOS (KP=4.00E-03 IS=3E-16 VTO=1)
.MODEL MI2 NMOS (KP=4.00E-03 IS=3E-16 VTO=0.9980)
.MODEL QOP PNP (BF=1.36E+02 IS=1E-14)
.MODEL QON NPN (BF=1.36E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
***********
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA01
* BEGIN OPAMP MACROMODEL PA16
* PINOUT ORDER +IN -IN RCL+ RCLC RCL- OUT +V -V
*                1   2  29   31   30   3   4  5
.SUBCKT PA16 1 2 29 31 30 3 4 5
* POSITIVE CURRENT LIMIT RESISTOR GOES FROM RCL+ TO RCLC
* NEGATIVE CURRENT LIMIT RESISTOR GOES FROM RCL- TO RCLC
* NOTE THAT CURRENT LIMIT RESISTORS DO NOT CONNECT TO THE SUPPLIES
* LIKE THEY DO IN THE PHYSICAL PART
J1 10 1 8 JI1
J2 11 2 9 JI2
R3 12 8 1.52E+03
R4 12 9 1.52E+03
I2 12 5 1.00E-04
C1 12 5 5.56E-13
R5 12 5 4.00E+06
R1 4 10 1.77E+03
R2 4 11 1.77E+03
C2 10 11 9.00E-12
I1 4 5 1.74E-02
G1 6 15 11 10 5.65E-04
G2 6 15 12 15 1.79E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 5.00E-12
G3 15 7 15 6 2.50E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 1.20E+00
D4 17 7 DD
V2 17 19 1.20E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 3.12E-11
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 1.19E-01
R13 22 24 1.19E-01
D5 23 25 DL
D6 26 24 DL
R9 27 29 1E3
R10 28 30 100
I3 18 23 9.47E-03
I4 24 19 9.47E-03
R15 31 3 4.18E-01
DC1 3 4 DO
DC2 5 3 DO
.MODEL DO D(CJO=10PF IS=5.25E-14 RS=5.71E-02)
RS1 29 31 1E6
RS2 30 31 1E6
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL JI1 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1)
.MODEL JI2 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1.0050)
.MODEL QOP PNP (BF=5.54E+02 IS=1E-14)
.MODEL QON NPN (BF=5.54E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
***********
* BEGIN OPAMP MACROMODEL PA162
* REVISION 1 28-AUGUST-2006 INITIAL RELEASE
* SYM=PA21
* PINOUT ORDER +IN -IN OUT +V -V
*                1  2   3   4  5
.SUBCKT PA162 1 2 3 4 5 
R4 9 12 7.39E+3 
R3 8 12 7.39E+3 
R1 4 10 8.85E+3 
R2 4 11 8.85E+3 
R5 12 5 111E6   
R6 6 0 100E+3   
R7 7 0 1000     
I2 12 5 16.6E-6 
C1 12 5 2.73E-12
C2 10 11 1E-12  
G1 6 0 11 10 113E-6     
G2 6 0 12 0 6.36E-9     
G3 0 7 0 6 25   
D1 6 0 DD       
D2 0 6 DD       
C3 6 7 4.4E-12  
I1 5 4 10.8E-3  
D3 7 16 DD      
D4 17 7 DD      
V1 18 16 1.63   
V2 17 19 1.63   
I3 4 23 6.3E-3  
I4 24 5 6.3E-3  
Q5 4 23 29 QON  
Q4 4 20 22 QON  
Q6 5 24 30 QOP  
Q3 5 20 21 QOP  
R58 51 20 50    
R8 7 50 50      
C54 20 0 .34E-9 
C4 50 0 .3E-9   
R15 31 3 .76    
E6 18 0 4 0 1   
E7 19 0 5 0 1   
E50 51 0 50 0 1 
Q1 10 1 8 QI1   
Q2 11 2 9 QI2   
Q8 26 28 31 QLP 
Q7 25 27 31 QLN 
D5 25 23 DL     
D6 24 26 DL     
R11 23 21 .26   
R13 22 24 .26   
RCLP 29 31 .26  
RCLN 31 30 .26  
R9 27 29 1000   
R10 28 30 1000
.MODEL DD D(CJO=0.1PF IS=1E-17) 
.MODEL DL D(CJO=3PF IS=1E-13)   
.MODEL QI1 NPN (BF=7.37E-01 IS=8E-16)   
.MODEL QI2 NPN (BF=6.67E-01 IS=8.45E-16)
.MODEL QOP PNP (BF=3.92E+02 IS=1E-14)   
.MODEL QON NPN (BF=3.92E+02 IS=1E-14)   
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
*************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA19
* BEGIN OPAMP MACROMODEL PA19
* PINOUT ORDER +IN -IN OUT +V -V COMP COMP PL ILC NL
*                1   2  3   4  5   6    7  29  31 30
.SUBCKT PA19 1 2 3 4 5 6 7 29 31 30
* THE COMPENSATION NETWORK IS CONNECTED FROM COMP TO COMP RATHER THAN FROM COMP TO OUT
* THE EXTERNAL POSITVE CURRENT LIMIT RESISTOR CONNECTS FROM PL TO ILC
* AND THE EXTERNAL NEGATIVE CURRENT LIMIT RESISTOR CONNECTS FROM NL TO ILC
*THEREFOR THE CURRENT LIMIT RESISTORS DO NOT CONNECT TO THE RAILS
*
M1 10 1 8 8 MI1
M2 11 2 9 9 MI2
R3 12 8 5.24E+01
R4 12 9 5.24E+01
I2 12 5 1.20E-02
C1 12 5 6.32E-13
R5 12 5 6.67E+04
R1 4 10 9.48E+01
R2 4 11 9.48E+01
C2 10 11 4.20E-11
I1 4 5 7.85E-02
G1 6 15 11 10 1.06E-02
G2 6 15 12 15 3.34E-07
R6 6 15 1.80E+04
D1 6 34 DD
D7 34 15 DD
D2 35 6 DD
D8 15 35 DD
C3 6 7 5.00E-12
G3 15 7 15 6 5.27E-02
R7 7 15 1E3
D3 7 16 DD
V1 18 16 9.50E-01
D4 17 7 DD
V2 17 19 9.50E-01
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 2.71E-11
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 1.19E-01
RCLP 29 31 1.19
RCLN 30 31 1.19
R13 22 24 1.19E-01
D5 23 25 DL
D6 26 24 DL
R9 27 29 1E3
R10 28 30 1E3
I3 18 23 9.47E-03
I4 24 19 9.47E-03
R15 31 3 8.72E-01
DC1 3 4 DO
DC2 5 3 DO
.MODEL DO D(CJO=10PF IS=5.25E-14 RS=5.71E-02)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MI1 NMOS (KP=2.36E-02 IS=3E-16 VTO=1)
.MODEL MI2 NMOS (KP=2.36E-02 IS=3E-16 VTO=0.9985)
.MODEL QOP PNP (BF=5.54E+02 IS=1E-14)
.MODEL QON NPN (BF=5.54E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-12)
.MODEL QLP PNP (BF=100 IS=1E-12)
* END OF OPAMP MACROMODEL
.ENDS
********************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA21
* BEGIN OPAMP MACROMODEL PA21
* PINOUT ORDER +IN -IN OUT +V -V
*                1  2   3   4  5
.SUBCKT PA21 1 2 3 4 5 
Q1 10 1 8 QI1
Q2 11 2 9 QI2
R3 12 8 7.39E+03
R4 12 9 7.39E+03
I2 12 5 3.61E-05
C1 12 5 2.73E-12
R5 12 5 1.11E+08
R1 4 10 8.85E+03
R2 4 11 8.85E+03
C2 10 11 9.00E-12
I1 4 5 3.70E-02
G1 6 15 11 10 1.13E-04
G2 6 15 12 15 6.36E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 3.00E-11
G3 15 7 15 6 8.85E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 1.60E+00
D4 17 7 DD
V2 17 19 1.60E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 3.08E-09
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 1.70E-01
RCLP 29 31 1.70E-01
RCLN 30 31 1.70E-01
R13 22 24 1.70E-01
D5 23 25 DL
D6 26 24 DL
R9 27 29 1E3
R10 28 30 1E3
I3 18 23 7.92E-03
I4 24 19 7.92E-03
R15 31 3 5.42E-01
RSN 3 34 1
CSN 34 5 0.1E-6
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL QI1 NPN (BF=6.55E+02 IS=8E-16)
.MODEL QI2 NPN (BF=4.24E+02 IS=8.46E-16)
.MODEL QOP PNP (BF=4.64E+02 IS=1E-14)
.MODEL QON NPN (BF=4.64E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
******************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA21
* BEGIN OPAMP MACROMODEL PA25
* PINOUT ORDER +IN -IN OUT +V -V
*                1   2  3   4  5
.SUBCKT PA25 1 2 3 4 5
Q1 10 1 8 QI1
Q2 11 2 9 QI2
R3 12 8 7.39E+03
R4 12 9 7.39E+03
I2 12 5 3.61E-05
C1 12 5 2.73E-12
R5 12 5 1.11E+08
R1 4 10 8.85E+03
R2 4 11 8.85E+03
C2 10 11 9.00E-12
I1 4 5 3.70E-02
G1 6 15 11 10 1.13E-04
G2 6 15 12 15 6.36E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 3.00E-11
G3 15 7 15 6 8.85E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 1.60E+00
D4 17 7 DD
V2 17 19 1.60E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 3.08E-09
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 1.70E-01
RCLP 29 31 1.70E-01
RCLN 30 31 1.70E-01
R13 22 24 1.70E-01
D5 23 25 DL
D6 26 24 DL
R9 27 29 1E3
R10 28 30 1E3
I3 18 23 7.92E-03
I4 24 19 7.92E-03
R15 31 3 5.42E-01
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL QI1 NPN (BF=6.55E+02 IS=8E-16)
.MODEL QI2 NPN (BF=4.24E+02 IS=8.46E-16)
.MODEL QOP PNP (BF=4.64E+02 IS=1E-14)
.MODEL QON NPN (BF=4.64E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
*************
*REVISION 3 26-JUN-2002
*REVISED E2, V1, DELETED V3 STOP G3 CURRENT GOING OUT THE +VS PIN.
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA26
* BEGIN OPAMP MACROMODEL PA26
* PINOUT ORDER +IN -IN OUT +V -V +VB ISEN
*                1   2  3   4  5  50  51
.SUBCKT PA26 1 2 3 4 5 50 51
Q1 10 1 8 QI1
Q2 11 2 9 QI2
R3 12 8 7.39E+03
R4 12 9 7.39E+03
I2 12 5 3.61E-05
C1 12 5 2.73E-12
R5 12 5 1.11E+08
R1 4 10 8.85E+03
R2 4 11 8.85E+03
C2 10 11 9.00E-12
I1 4 5 2.50E-02
G1 6 15 11 10 1.13E-04
G2 6 15 12 15 6.36E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 3.00E-11
G3 15 7 15 6 8.85E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 1.10E+00
D4 17 7 DD
V2 17 19 1.60E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 3.08E-09
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 51 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 1.70E-01
RCLP 29 31 1.70E-01
RCLN 30 31 1.70E-01
R13 22 24 1.70E-01
D5 23 25 DL
D6 26 24 DL
R9 27 29 1E3
R10 28 30 1E3
I3 18 23 7.92E-03
I4 24 19 7.92E-03
R15 31 3 5.42E-01
E4 54 18 50 4 .15
V4 54 53 1.6
D8 7 53 DD
I5 50 5 12E-03
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL QI1 NPN (BF=6.55E+02 IS=8E-16)
.MODEL QI2 NPN (BF=4.24E+02 IS=8.46E-16)
.MODEL QOP PNP (BF=4.64E+02 IS=1E-14)
.MODEL QON NPN (BF=4.64E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA04
* BEGIN OPAMP MACROMODEL PA33
* PINOUT ORDER  +IN -IN OUT ILIM-10 ILIM-11 +VB -VB
* PINOUT ORDER CONTINUED  COMP COMP +VS -VS
.SUBCKT PA33 1 2 3 33 31 4 5 6 7 36 37
M1 10 1 8 8 MI1
M2 11 2 9 9 MI2
R3 12 8 5.40E+01
R4 12 9 5.40E+01
I2 12 5 8.99E-03
C1 12 5 1.76E-12
R5 12 5 2.76E+06
R1 4 10 1.26E+02
R2 4 11 1.26E+02
C2 10 11 2.10E-10
I1 4 5 3.69E-02
G1 6 15 11 10 7.91E-03
G2 6 15 12 15 7.91E-08
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 5.00E-12
G3 15 7 15 6 1.59E-01
R7 7 15 1E3
D3 7 16 DD
V1 18 16 6.70E+00
D4 17 7 DD
V2 17 19 6.70E+00
RE1 15 0 0.001
E2 38 0 4 0 1
E3 39 0 5 0 1
R8 7 20 50
C4 20 15 3.79E-10
Q3 37 20 21 QOP
Q4 36 20 22 QON
Q5 36 21 29 QON
Q6 37 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 31 1E3
R10 28 31 1E3
E4 41 36 38 36 1
E5 42 37 39 37 1
E6 18 0 41 0 1
E7 19 0 42 0 1
RY1 38 0 10E6
RY2 39 0 10E6
RY3 41 0 10E6
RY4 42 0 10E6
I3 36 21 7.15E-03
I4 22 37 7.15E-03
R15 29 3 1.58E-01
DC1 29 36 DO
DC2 37 29 DO
I5 36 37 2.25E-02
.MODEL DO D(CJO=10PF IS=3.99E-13 RS=7.52E-03)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MI1 NMOS (KP=1.38E-02 IS=3E-16 VTO=1)
.MODEL MI2 NMOS (KP=1.38E-02 IS=3E-16 VTO=0.9950)
.MODEL QOP PNP (BF=5.58E+03 IS=1E-14)
.MODEL QON NPN (BF=5.58E+03 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
*************
*REVISION 3 26-JUN-2002
*REVISED E2, V1, DELETED V3 STOP G3 CURRENT GOING OUT THE +VS PIN.
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA26
* BEGIN OPAMP MACROMODEL PA34
* PINOUT ORDER +IN -IN OUT +V -V +VB ISEN
*                1   2  3   4  5  50  51
.SUBCKT PA34 1 2 3 4 5 50 51
Q1 10 1 8 QI1
Q2 11 2 9 QI2
R3 12 8 7.39E+03
R4 12 9 7.39E+03
I2 12 5 3.61E-05
C1 12 5 2.73E-12
R5 12 5 1.11E+08
R1 4 10 8.85E+03
R2 4 11 8.85E+03
C2 10 11 9.00E-12
I1 4 5 2.50E-02
G1 6 15 11 10 1.13E-04
G2 6 15 12 15 6.36E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 3.00E-11
G3 15 7 15 6 8.85E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 1.10E+00
D4 17 7 DD
V2 17 19 1.60E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 3.08E-09
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 51 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 1.70E-01
RCLP 29 31 1.70E-01
RCLN 30 31 1.70E-01
R13 22 24 1.70E-01
D5 23 25 DL
D6 26 24 DL
R9 27 29 1E3
R10 28 30 1E3
I3 18 23 7.92E-03
I4 24 19 7.92E-03
R15 31 3 5.42E-01
E4 54 18 50 4 .15
V4 54 53 1.6
D8 7 53 DD
I5 50 5 12E-03
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL QI1 NPN (BF=6.55E+02 IS=8E-16)
.MODEL QI2 NPN (BF=4.24E+02 IS=8.46E-16)
.MODEL QOP PNP (BF=4.64E+02 IS=1E-14)
.MODEL QON NPN (BF=4.64E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
******************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA21
* BEGIN OPAMP MACROMODEL PA35AMP
* PINOUT ORDER +IN -IN OUT +V -V
*                1   2  3   4  5
.SUBCKT PA35AMP 1 2 3 4 5
Q1 10 1 8 QI1
Q2 11 2 9 QI2
R3 12 8 7.39E+03
R4 12 9 7.39E+03
I2 12 5 3.61E-05
C1 12 5 2.73E-12
R5 12 5 1.11E+08
R1 4 10 8.85E+03
R2 4 11 8.85E+03
C2 10 11 9.00E-12
I1 4 5 3.70E-02
G1 6 15 11 10 1.13E-04
G2 6 15 12 15 6.36E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 3.00E-11
G3 15 7 15 6 8.85E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 1.60E+00
D4 17 7 DD
V2 17 19 1.60E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 3.08E-09
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 1.70E-01
RCLP 29 31 1.70E-01
RCLN 30 31 1.70E-01
R13 22 24 1.70E-01
D5 23 25 DL
D6 26 24 DL
R9 27 29 1E3
R10 28 30 1E3
I3 18 23 7.92E-03
I4 24 19 7.92E-03
R15 31 3 5.42E-01
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL QI1 NPN (BF=6.55E+02 IS=8E-16)
.MODEL QI2 NPN (BF=4.24E+02 IS=8.46E-16)
.MODEL QOP PNP (BF=4.64E+02 IS=1E-14)
.MODEL QON NPN (BF=4.64E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
*************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
* BEGIN OPAMP MACROMODEL PA35BUF
* PINOUT ORDER +IN OUT +V -V
*                1  3   4  5
.SUBCKT PA35BUF 1 3 4 5
Q1 10 1 8 QI1
Q2 11 3 9 QI2
R3 12 8 7.39E+03
R4 12 9 7.39E+03
I2 12 5 3.61E-05
C1 12 5 2.73E-12
R5 12 5 1.11E+08
R1 4 10 8.85E+03
R2 4 11 8.85E+03
C2 10 11 9.00E-12
I1 4 5 3.70E-02
G1 6 15 11 10 1.13E-04
G2 6 15 12 15 6.36E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 3.00E-11
G3 15 7 15 6 8.85E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 1.60E+00
D4 17 7 DD
V2 17 19 1.60E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 3.08E-09
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 1.70E-01
RCLP 29 31 1.70E-01
RCLN 30 31 1.70E-01
R13 22 24 1.70E-01
D5 23 25 DL
D6 26 24 DL
R9 27 29 1E3
R10 28 30 1E3
I3 18 23 7.92E-03
I4 24 19 7.92E-03
R15 31 3 5.42E-01
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL QI1 NPN (BF=6.55E+02 IS=8E-16)
.MODEL QI2 NPN (BF=4.24E+02 IS=8.46E-16)
.MODEL QOP PNP (BF=4.64E+02 IS=1E-14)
.MODEL QON NPN (BF=4.64E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
*************
*REVISION 3 26-JUN-2002
*REVISED E2, V1, DELETED V3 STOP G3 CURRENT GOING OUT THE +VS PIN.
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA26
* BEGIN OPAMP MACROMODEL PA37
* PINOUT ORDER +IN -IN OUT +V -V +VB ISEN
*                1   2  3   4  5  50  51
.SUBCKT PA37 1 2 3 4 5 50 51
Q1 10 1 8 QI1
Q2 11 2 9 QI2
R3 12 8 7.39E+03
R4 12 9 7.39E+03
I2 12 5 3.61E-05
C1 12 5 2.73E-12
R5 12 5 1.11E+08
R1 4 10 8.85E+03
R2 4 11 8.85E+03
C2 10 11 9.00E-12
I1 4 5 2.50E-02
G1 6 15 11 10 1.13E-04
G2 6 15 12 15 6.36E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 3.00E-11
G3 15 7 15 6 8.85E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 1.10E+00
D4 17 7 DD
V2 17 19 1.60E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 3.08E-09
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 51 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 1.70E-01
RCLP 29 31 1.70E-01
RCLN 30 31 1.70E-01
R13 22 24 1.70E-01
D5 23 25 DL
D6 26 24 DL
R9 27 29 1E3
R10 28 30 1E3
I3 18 23 7.92E-03
I4 24 19 7.92E-03
R15 31 3 5.42E-01
E4 54 18 50 4 .15
V4 54 53 1.6
D8 7 53 DD
I5 50 5 12E-03
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL QI1 NPN (BF=6.55E+02 IS=8E-16)
.MODEL QI2 NPN (BF=4.24E+02 IS=8.46E-16)
.MODEL QOP PNP (BF=4.64E+02 IS=1E-14)
.MODEL QON NPN (BF=4.64E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
*************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA09
* BEGIN OPAMP MACROMODEL PA40
* PINOUT ORDER +IN -IN OUT +V -V COMP COMP
*                1   2  3   4  5   6    7
.SUBCKT PA40 1 2 3 4 5 6 7
M1 10 1 8 8 MI1
M2 11 2 9 9 MI2
R3 12 8 2.95E+03
R4 12 9 2.95E+03
I2 12 5 2.90E-04
C1 12 5 7.78E-13
R5 12 5 1.38E+07
R1 4 10 3.20E+03
R2 4 11 3.20E+03
C2 10 11 1.66E-11
I1 4 5 -8.81E-05
G1 6 15 11 10 3.13E-04
G2 6 15 12 15 5.56E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 5.00E-12
G3 15 7 15 6 5.69E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 3.20E+00
D4 17 7 DD
V2 17 19 6.70E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 9.35E-11
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
M3 25 27 3 3 MLN
M4 26 28 3 3 MLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 1.20E-03
I4 22 19 1.20E-03
R15 29 3 7.50E+01
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=8.40E-16 RS=3.57E+00)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MI1 NMOS (KP=4.00E-03 IS=3E-16 VTO=1)
.MODEL MI2 NMOS (KP=4.00E-03 IS=3E-16 VTO=0.9850)
.MODEL MLN NMOS (KP=5.00E-03 IS=3E-16 VTO=2.5)
.MODEL MLP PMOS (KP=5.00E-03 IS=3E-16 VTO=-2.5)
.MODEL QOP PNP (BF=7.01E+01 IS=1E-14)
.MODEL QON NPN (BF=7.01E+01 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.*SYM=PA85
* BEGIN OPAMP MACROMODEL PA41
* PINOUT ORDER +IN -IN CL OUT +V -V COMP COMP
*                1   2  3  33  4  5   6    7
.SUBCKT PA41 1 2 3 33 4 5 6 7
M1 10 1 8 8 MI1
M2 11 2 9 9 MI2
R3 12 8 2.95E+03
R4 12 9 2.95E+03
I2 12 5 2.90E-04
C1 12 5 7.78E-13
R5 12 5 1.38E+07
R1 4 10 3.20E+03
R2 4 11 3.20E+03
C2 10 11 1.66E-11
I1 4 5 -8.81E-05
G1 6 15 11 10 3.13E-04
G2 6 15 12 15 5.56E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 5.00E-12
G3 15 7 15 6 5.69E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 3.20E+00
D4 17 7 DD
V2 17 19 6.70E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 9.35E-11
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
M3 25 27 33 33 MLN
M4 26 28 33 33 MLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 1.20E-03
I4 22 19 1.20E-03
R15 29 3 7.50E+01
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=8.40E-16 RS=3.57E+00)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MI1 NMOS (KP=4.00E-03 IS=3E-16 VTO=1)
.MODEL MI2 NMOS (KP=4.00E-03 IS=3E-16 VTO=0.9850)
.MODEL MLN NMOS (KP=5.00E-03 IS=3E-16 VTO=2.5)
.MODEL MLP PMOS (KP=5.00E-03 IS=3E-16 VTO=-2.5)
.MODEL QOP PNP (BF=7.01E+01 IS=1E-14)
.MODEL QON NPN (BF=7.01E+01 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
*************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA85
* BEGIN OPAMP MACROMODEL PA42
* PINOUT ORDER +IN -IN CL OUT +V -V COMP COMP
*                1   2  3  33  4  5   6    7
.SUBCKT PA42 1 2 3 33 4 5 6 7
M1 10 1 8 8 MI1
M2 11 2 9 9 MI2
R3 12 8 2.95E+03
R4 12 9 2.95E+03
I2 12 5 2.90E-04
C1 12 5 7.78E-13
R5 12 5 1.38E+07
R1 4 10 3.20E+03
R2 4 11 3.20E+03
C2 10 11 1.66E-11
I1 4 5 -8.81E-05
G1 6 15 11 10 3.13E-04
G2 6 15 12 15 5.56E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 5.00E-12
G3 15 7 15 6 5.69E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 3.20E+00
D4 17 7 DD
V2 17 19 6.70E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 9.35E-11
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
M3 25 27 33 33 MLN
M4 26 28 33 33 MLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 1.20E-03
I4 22 19 1.20E-03
R15 29 3 7.50E+01
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=8.40E-16 RS=3.57E+00)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MI1 NMOS (KP=4.00E-03 IS=3E-16 VTO=1)
.MODEL MI2 NMOS (KP=4.00E-03 IS=3E-16 VTO=0.9850)
.MODEL MLN NMOS (KP=5.00E-03 IS=3E-16 VTO=2.5)
.MODEL MLP PMOS (KP=5.00E-03 IS=3E-16 VTO=-2.5)
.MODEL QOP PNP (BF=7.01E+01 IS=1E-14)
.MODEL QON NPN (BF=7.01E+01 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
*************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA85
* BEGIN OPAMP MACROMODEL PA44
* PINOUT ORDER +IN -IN CL OUT +V -V COMP COMP
*                1   2  3  33  4  5   6    7
.SUBCKT PA44 1 2 3 33 4 5 6 7
M1 10 1 8 8 MI1
M2 11 2 9 9 MI2
R3 12 8 2.95E+03
R4 12 9 2.95E+03
I2 12 5 2.90E-04
C1 12 5 7.78E-13
R5 12 5 1.38E+07
R1 4 10 3.20E+03
R2 4 11 3.20E+03
C2 10 11 1.66E-11
I1 4 5 -8.81E-05
G1 6 15 11 10 3.13E-04
G2 6 15 12 15 5.56E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 5.00E-12
G3 15 7 15 6 5.69E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 3.20E+00
D4 17 7 DD
V2 17 19 6.70E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 9.35E-11
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
M3 25 27 33 33 MLN
M4 26 28 33 33 MLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 1.20E-03
I4 22 19 1.20E-03
R15 29 3 7.50E+01
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=8.40E-16 RS=3.57E+00)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MI1 NMOS (KP=4.00E-03 IS=3E-16 VTO=1)
.MODEL MI2 NMOS (KP=4.00E-03 IS=3E-16 VTO=0.9850)
.MODEL MLN NMOS (KP=5.00E-03 IS=3E-16 VTO=2.5)
.MODEL MLP PMOS (KP=5.00E-03 IS=3E-16 VTO=-2.5)
.MODEL QOP PNP (BF=7.01E+01 IS=1E-14)
.MODEL QON NPN (BF=7.01E+01 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
***********
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
* BEGIN OPAMP MACROMODEL PA50
* PINOUT ORDER  +IN -IN OUT +VB -VB +VS -VS
.SUBCKT PA50 1 2 3 4 5 36 37
J1 10 1 8 JI1
J2 11 2 9 JI2
R3 12 8 1.34E+03
R4 12 9 1.34E+03
I2 12 5 4.50E-04
C1 12 5 5.00E-13
R5 12 5 5.45E+06
R1 4 10 1.59E+03
R2 4 11 1.59E+03
C2 10 11 1.67E-11
I1 4 5 2.64E-02
G1 6 15 11 10 6.28E-04
G2 6 15 12 15 2.81E-08
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 7.50E-12
G3 15 7 15 6 1.00E+01
R7 7 15 1E3
D3 7 16 DD
V1 18 16 5.50E+00
D4 17 7 DD
V2 17 19 5.50E+00
RE1 15 0 0.001
E2 38 0 4 0 1
E3 39 0 5 0 1
R8 7 20 50
C4 20 15 5.80E-11
Q3 37 20 21 QOP
Q4 36 20 22 QON
Q5 36 21 29 QON
Q6 37 22 29 QOP
E4 41 36 38 36 0.69
E5 42 37 39 37 0.69
E6 18 0 41 0 1
E7 19 0 42 0 1
RY1 38 0 10E6
RY2 39 0 10E6
RY3 41 0 10E6
RY4 42 0 10E6
I3 36 21 5.36E-03
I4 22 37 5.36E-03
I5 37 36 1.0E-02
R15 29 3 8.5E-02
DC1 29 36 DO
DC2 37 29 DO
.MODEL DO D(CJO=10PF IS=1.26E-12 RS=2.38E-03)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL JI1 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1)
.MODEL JI2 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1.0050)
.MODEL QOP PNP (BF=2.35E+04 IS=1E-14)
.MODEL QON NPN (BF=2.35E+04 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
************
*REVISION 3 12-3-2004
*CHANGED FROM CLASS AB TO CLASS C OPERATION
*REVISED CURRENT LIMIT TO MAKE SYMMETRIC
*REMOVED RE1
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA01
* BEGIN OPAMP MACROMODEL PA51
* PINOUT ORDER +IN -IN RCL+ RCLC RCL- OUT +V -V
*               1   2   29   31   30   3   4  5
.SUBCKT PA51 1 2 29 31 30 3 4 5
* POSITIVE CURRENT LIMIT RESISTOR GOES FROM RCL+ TO RCLC
* NEGATIVE CURRENT LIMIT RESISTOR GOES FROM RCL- TO RCLC
* NOTE THAT CURRENT LIMIT RESISTORS DO NOT CONNECT TO THE OUTPUT
* LIKE THEY DO IN THE PHYSICAL PART
* JUST LIKE THE REAL CLASS C PART SMALL SIGNAL ANALYSIS WILL APPEAR 
* TO HAVE SIGNIFICANTLY LOW GAIN UNLESS THE OUTPUT IS LOADED SUCH
* THAT OUTPUT STAGE CURRENT NEVER CHANGES POLARITY
Q1 10 1 8 QI1
Q2 11 2 9 QI2
R3 12 8 2.71E+03
R4 12 9 2.71E+03
I2 12 5 5.72E-05
C1 12 5 4.00E-12
R5 12 5 1.57E+08
R1 4 10 3.62E+03
R2 4 11 3.62E+03
C2 10 11 1.10E-11
I1 4 5 3E-03
G1 6 0 11 10 2.76E-04
G2 6 0 12 0 2.76E-09
R6 6 0 1.00E+05
D1 6 0 DD
D2 0 6 DD
C3 6 7 2.20E-11
G3 0 7 0 6 4.06E+00
R7 7 0 1E3
D3 7 16 DD
V1 18 16 3.95E+00
D4 17 7 DD
V2 17 19 3.15E+00
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 0 3.60E-10
Q3 19 20 71 QOP
Q4 18 20 72 QON
V3 71 21 .65
V4 22 72 .65
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 5.41E-02
R13 22 24 5.41E-02
D5 23 25 DL
D6 26 24 DL
R9 27 29 280
R10 28 30 280
I3 18 23 1.40E-02
I4 24 19 1.40E-02
R15 31 3 1.25E-01
DC1 3 4 DO
DC2 5 3 DO
.MODEL DO D(CJO=10PF IS=1.15E-13 RS=2.60E-02)
RS1 29 31 1E6
RS2 30 31 1E6
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL QI1 NPN (BF=1.91E+03 IS=8E-16)
.MODEL QI2 NPN (BF=1.90E+03 IS=8.62E-16)
.MODEL QOP PNP (BF=8.22E+02 IS=1E-14)
.MODEL QON NPN (BF=8.22E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-12)
.MODEL QLP PNP (BF=100 IS=1E-12)
* END OF OPAMP MACROMODEL
.ENDS
**********
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
* BEGIN OPAMP MACROMODEL PA52
* PINOUT ORDER  +IN -IN OUT +VB -VB +VS -VS
.SUBCKT PA52 1 2 3 4 5 36 37
J1 10 1 8 JI1
J2 11 2 9 JI2
R3 12 8 1.34E+03
R4 12 9 1.34E+03
I2 12 5 3.30E-04
C1 12 5 5.00E-13
R5 12 5 1.09E+07
R1 4 10 1.59E+03
R2 4 11 1.59E+03
C2 10 11 2.2E-11
I1 4 5 2.64E-02
G1 6 15 11 10 6.28E-04
G2 6 15 12 15 1.99E-08
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 5.5E-12
G3 15 7 15 6 1.00E+01
R7 7 15 1E3
D3 7 16 DD
V1 18 16 5.50E+00
D4 17 7 DD
V2 17 19 5.50E+00
RE1 15 0 0.001
E2 38 0 4 0 1
E3 39 0 5 0 1
R8 7 20 50
C4 20 15 3.80E-11
Q3 37 20 21 QOP
Q4 36 20 22 QON
Q5 36 21 29 QON
Q6 37 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 31 1E3
R10 28 31 1E3
E4 41 36 38 36 0.69
E5 42 37 39 37 0.69
E6 18 0 41 0 1
E7 19 0 42 0 1
RY1 38 0 10E6
RY2 39 0 10E6
RY3 41 0 10E6
RY4 42 0 10E6
I3 36 21 5.36E-03
I4 22 37 5.36E-03
I5 37 36 1.0E-02
R15 29 3 8.50E-02
DC1 29 36 DO
DC2 37 29 DO
.MODEL DO D(CJO=10PF IS=1.05E-12 RS=2.86E-03)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL JI1 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1)
.MODEL JI2 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1.0050)
.MODEL QOP PNP (BF=1.96E+04 IS=1E-14)
.MODEL QON NPN (BF=1.96E+04 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
*************
* BEGIN OPAMP MACROMODEL PA60
* REVISION 1 3-MARCH-2004 INITIAL RELEASE
* SYM=PA21
* PINOUT ORDER +IN -IN OUT +V -V
*                1  2   3   4  5
.SUBCKT PA60 1 2 3 4 5 
R4 9 12 7.39E+3 
R3 8 12 7.39E+3 
R1 4 10 8.85E+3 
R2 4 11 8.85E+3 
R5 12 5 111E6   
R6 6 0 100E+3   
R7 7 0 1000     
I2 12 5 16.6E-6 
C1 12 5 2.73E-12
C2 10 11 1E-12  
G1 6 0 11 10 113E-6     
G2 6 0 12 0 6.36E-9     
G3 0 7 0 6 25   
D1 6 0 DD       
D2 0 6 DD       
C3 6 7 4.4E-12  
I1 5 4 10.8E-3  
D3 7 16 DD      
D4 17 7 DD      
V1 18 16 1.63   
V2 17 19 1.63   
I3 4 23 6.3E-3  
I4 24 5 6.3E-3  
Q5 4 23 29 QON  
Q4 4 20 22 QON  
Q6 5 24 30 QOP  
Q3 5 20 21 QOP  
R58 51 20 50    
R8 7 50 50      
C54 20 0 .34E-9 
C4 50 0 .3E-9   
R15 31 3 .76    
E6 18 0 4 0 1   
E7 19 0 5 0 1   
E50 51 0 50 0 1 
Q1 10 1 8 QI1   
Q2 11 2 9 QI2   
Q8 26 28 31 QLP 
Q7 25 27 31 QLN 
D5 25 23 DL     
D6 24 26 DL     
R11 23 21 .26   
R13 22 24 .26   
RCLP 29 31 .26  
RCLN 31 30 .26  
R9 27 29 1000   
R10 28 30 1000
.MODEL DD D(CJO=0.1PF IS=1E-17) 
.MODEL DL D(CJO=3PF IS=1E-13)   
.MODEL QI1 NPN (BF=7.37E-01 IS=8E-16)   
.MODEL QI2 NPN (BF=6.67E-01 IS=8.45E-16)
.MODEL QOP PNP (BF=3.92E+02 IS=1E-14)   
.MODEL QON NPN (BF=3.92E+02 IS=1E-14)   
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
***********
*REVISION 1 12-3-2004
*INITIAL RELEASE COPIED FROM PA51 REVISION 3
*SYM=PA01
* BEGIN OPAMP MACROMODEL PA61
* PINOUT ORDER +IN -IN RCL+ RCLC RCL- OUT +V -V
*               1   2   29   31   30   3   4  5
.SUBCKT PA61 1 2 29 31 30 3 4 5
* POSITIVE CURRENT LIMIT RESISTOR GOES FROM RCL+ TO RCLC
* NEGATIVE CURRENT LIMIT RESISTOR GOES FROM RCL- TO RCLC
* NOTE THAT CURRENT LIMIT RESISTORS DO NOT CONNECT TO THE OUTPUT
* LIKE THEY DO IN THE PHYSICAL PART
* JUST LIKE THE REAL CLASS C PART SMALL SIGNAL ANALYSIS WILL APPEAR 
* TO HAVE SIGNIFICANTLY LOW GAIN UNLESS THE OUTPUT IS LOADED SUCH
* THAT OUTPUT STAGE CURRENT NEVER CHANGES POLARITY
Q1 10 1 8 QI1
Q2 11 2 9 QI2
R3 12 8 2.71E+03
R4 12 9 2.71E+03
I2 12 5 5.72E-05
C1 12 5 4.00E-12
R5 12 5 1.57E+08
R1 4 10 3.62E+03
R2 4 11 3.62E+03
C2 10 11 1.10E-11
I1 4 5 3E-03
G1 6 0 11 10 2.76E-04
G2 6 0 12 0 2.76E-09
R6 6 0 1.00E+05
D1 6 0 DD
D2 0 6 DD
C3 6 7 2.20E-11
G3 0 7 0 6 4.06E+00
R7 7 0 1E3
D3 7 16 DD
V1 18 16 3.95E+00
D4 17 7 DD
V2 17 19 3.15E+00
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 0 3.60E-10
Q3 19 20 71 QOP
Q4 18 20 72 QON
V3 71 21 .65
V4 22 72 .65
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 5.41E-02
R13 22 24 5.41E-02
D5 23 25 DL
D6 26 24 DL
R9 27 29 280
R10 28 30 280
I3 18 23 1.40E-02
I4 24 19 1.40E-02
R15 31 3 1.25E-01
DC1 3 4 DO
DC2 5 3 DO
.MODEL DO D(CJO=10PF IS=1.15E-13 RS=2.60E-02)
RS1 29 31 1E6
RS2 30 31 1E6
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL QI1 NPN (BF=1.91E+03 IS=8E-16)
.MODEL QI2 NPN (BF=1.90E+03 IS=8.62E-16)
.MODEL QOP PNP (BF=8.22E+02 IS=1E-14)
.MODEL QON NPN (BF=8.22E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-12)
.MODEL QLP PNP (BF=100 IS=1E-12)
* END OF OPAMP MACROMODEL
.ENDS
*************
* BEGIN OPAMP MACROMODEL PA62
* REVISION 1 28-AUGUST-2006 INITIAL RELEASE
* SYM=PA21
* PINOUT ORDER +IN -IN OUT +V -V
*                1  2   3   4  5
.SUBCKT PA62 1 2 3 4 5 
R4 9 12 7.39E+3 
R3 8 12 7.39E+3 
R1 4 10 8.85E+3 
R2 4 11 8.85E+3 
R5 12 5 111E6   
R6 6 0 100E+3   
R7 7 0 1000     
I2 12 5 16.6E-6 
C1 12 5 2.73E-12
C2 10 11 1E-12  
G1 6 0 11 10 113E-6     
G2 6 0 12 0 6.36E-9     
G3 0 7 0 6 25   
D1 6 0 DD       
D2 0 6 DD       
C3 6 7 4.4E-12  
I1 5 4 10.8E-3  
D3 7 16 DD      
D4 17 7 DD      
V1 18 16 1.63   
V2 17 19 1.63   
I3 4 23 6.3E-3  
I4 24 5 6.3E-3  
Q5 4 23 29 QON  
Q4 4 20 22 QON  
Q6 5 24 30 QOP  
Q3 5 20 21 QOP  
R58 51 20 50    
R8 7 50 50      
C54 20 0 .34E-9 
C4 50 0 .3E-9   
R15 31 3 .76    
E6 18 0 4 0 1   
E7 19 0 5 0 1   
E50 51 0 50 0 1 
Q1 10 1 8 QI1   
Q2 11 2 9 QI2   
Q8 26 28 31 QLP 
Q7 25 27 31 QLN 
D5 25 23 DL     
D6 24 26 DL     
R11 23 21 .26   
R13 22 24 .26   
RCLP 29 31 .26  
RCLN 31 30 .26  
R9 27 29 1000   
R10 28 30 1000
.MODEL DD D(CJO=0.1PF IS=1E-17) 
.MODEL DL D(CJO=3PF IS=1E-13)   
.MODEL QI1 NPN (BF=7.37E-01 IS=8E-16)   
.MODEL QI2 NPN (BF=6.67E-01 IS=8.45E-16)
.MODEL QOP PNP (BF=3.92E+02 IS=1E-14)   
.MODEL QON NPN (BF=3.92E+02 IS=1E-14)   
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
*************
*REVISION 2 26-NOV-2004
*REVISE GAIN AND PHASE TO MATCH NEW DATA SHEET
*MAKE ILIMIT SYMMETRIC
*REVISION 1 6-MAY-2004 INITIAL RELEASE
*SYM=PA01
* BEGIN OPAMP MACROMODEL PA73
* PINOUT ORDER +IN -IN RCL+ RCLC RCL- OUT +V -V
*                1   2  29   31   30   3   4  5
.SUBCKT PA73 1 2 29 31 30 3 4 5
* POSITIVE CURRENT LIMIT RESISTOR GOES FROM RCL+ TO RCLC
* NEGATIVE CURRENT LIMIT RESISTOR GOES FROM RCL- TO RCLC
* NOTE THAT CURRENT LIMIT RESISTORS DO NOT CONNECT TO THE OUTPUT
* LIKE THEY DO IN THE PHYSICAL PART
Q1 10 1 8 QI1
Q2 11 2 9 QI2
R3 12 8 2.68E+03
R4 12 9 2.68E+03
I2 12 5 31E-06
C1 12 5 1.43E-12
R5 12 5 2.5E+08
R1 4 10 3.98E+03
R2 4 11 3.98E+03
C2 10 11 5E-12
I1 4 5 2.6E-03
G1 6 0 11 10 2.51E-04
G2 6 0 12 0 1.41E-09
R6 6 0 1.00E+05
D1 6 0 DD
D2 0 6 DD
C3 6 7 10E-12
G3 0 7 0 6 4.5E+00
R7 7 0 1E3
D3 7 16 DD
V1 18 16 4.70E+00
D4 17 7 DD
V2 17 19 4.70E+00
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 0 278E-12
Q3 19 20 71 QOP
Q4 18 20 72 QON
V3 71 21 .65
V4 22 72 .65
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 1.08E-01
R13 22 24 1.08E-01
D5 23 25 DL
D6 26 24 DL
R9 27 29 550
R10 28 30 550
I3 18 23 9.93E-03
I4 24 19 9.93E-03
R15 31 3 6.67E-01
DC1 3 4 DO
DC2 5 3 DO
.MODEL DO D(CJO=10PF IS=5.77E-14 RS=5.19E-02)
RS1 29 31 1E6
RS2 30 31 1E6
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL QI1 NPN (BF=2.22E+03 IS=8E-16)
.MODEL QI2 NPN (BF=1.33E+03 IS=9.54E-16)
.MODEL QOP PNP (BF=5.82E+02 IS=1E-14)
.MODEL QON NPN (BF=5.82E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-12)
.MODEL QLP PNP (BF=100 IS=1E-12)
* END OF OPAMP MACROMODEL
.ENDS
***********
* BEGIN OPAMP MACROMODEL PA74
* REVISION 1 15-DECEMBER-2003 INITIAL RELEASE
* SYM=PA21
* PINOUT ORDER +IN -IN OUT +V -V
*                1  2   3   4  5
.SUBCKT PA74 1 2 3 4 5 
R4 9 12 7.39E+3 
R3 8 12 7.39E+3 
R1 4 10 8.85E+3 
R2 4 11 8.85E+3 
R5 12 5 111E6   
R6 6 0 100E+3   
R7 7 0 1000     
I2 12 5 16.6E-6 
C1 12 5 2.73E-12
C2 10 11 1E-12  
G1 6 0 11 10 113E-6     
G2 6 0 12 0 6.36E-9     
G3 0 7 0 6 25   
D1 6 0 DD       
D2 0 6 DD       
C3 6 7 4.4E-12  
I1 5 4 10.8E-3  
D3 7 16 DD      
D4 17 7 DD      
V1 18 16 1.63   
V2 17 19 1.63   
I3 4 23 6.3E-3  
I4 24 5 6.3E-3  
Q5 4 23 29 QON  
Q4 4 20 22 QON  
Q6 5 24 30 QOP  
Q3 5 20 21 QOP  
R58 51 20 50    
R8 7 50 50      
C54 20 0 .34E-9 
C4 50 0 .3E-9   
R15 31 303 .76    
E6 18 0 4 0 1   
E7 19 0 5 0 1   
E50 51 0 50 0 1 
Q1 10 1 8 QI1   
Q2 11 2 9 QI2   
Q8 26 52 31 QLP 
Q7 25 53 31 QLN 
D5 25 23 DL     
D6 24 26 DL     
R11 23 21 .26   
R13 22 24 .26   
RCLP 29 31 .26  
RCLN 31 30 .26  
R9 53 29 1000   
R10 52 30 1000
*BUFFER 1
R104 109 112 7.39E+3 
R103 108 112 7.39E+3 
R101 4 110 8.85E+3 
R102 4 111 8.85E+3 
R105 112 5 111E6   
R106 106 0 100E+3   
R107 107 0 1000     
I102 112 5 16.6E-6 
C101 112 5 2.73E-12
C102 110 111 1E-12  
G101 106 0 111 10 113E-6     
G102 106 0 112 0 6.36E-9     
G103 0 107 0 106 25   
D101 106 0 DD       
D102 0 106 DD       
C103 106 107 4.4E-12  
I101 5 4 10.8E-3  
D103 107 116 DD      
D104 117 107 DD      
V101 118 116 1.63   
V102 117 119 1.63   
I103 4 123 6.3E-3  
I104 124 5 6.3E-3  
Q105 4 123 129 QON  
Q104 4 120 122 QON  
Q106 5 124 130 QOP  
Q103 5 120 121 QOP  
R158 151 120 50    
R108 107 150 50      
C154 120 0 .34E-9 
C104 150 0 .3E-9   
R115 131 103 .76    
E106 118 0 4 0 1   
E107 119 0 5 0 1   
E150 151 0 150 0 1 
Q101 110 303 108 QI1   
Q102 111 103 109 QI2   
Q108 126 152 131 QLP 
Q107 125 153 131 QLN 
D105 125 123 DL     
D106 124 126 DL     
R111 123 121 .26   
R113 122 124 .26   
R1CLP 129 131 .26  
R1CLN 131 130 .26  
R109 153 129 1000   
R110 152 130 1000
*BUFFER2
R204 209 212 7.39E+3 
R203 208 212 7.39E+3 
R201 4 210 8.85E+3 
R202 4 211 8.85E+3 
R205 12 5 111E6   
R206 206 0 100E+3   
R207 207 0 1000     
I202 212 5 16.6E-6 
C201 212 5 2.73E-12
C202 210 211 1E-12  
G201 206 0 211 10 113E-6     
G202 206 0 212 0 6.36E-9     
G203 0 207 0 206 25   
D201 206 0 DD       
D202 0 206 DD       
C203 206 207 4.4E-12  
I201 5 4 10.8E-3  
D203 207 216 DD      
D204 217 207 DD      
V201 218 216 1.63   
V202 217 219 1.63   
I203 4 223 6.3E-3  
I204 224 5 6.3E-3  
Q205 4 223 229 QON  
Q204 4 220 222 QON  
Q206 5 224 230 QOP  
Q203 5 220 221 QOP  
R258 251 220 50    
R208 207 250 50      
C254 220 0 .34E-9 
C204 250 0 .3E-9   
R215 231 203 .76    
E206 218 0 4 0 1   
E207 219 0 5 0 1   
E250 251 0 250 0 1 
Q201 210 303 208 QI1   
Q202 211 203 209 QI2   
Q208 226 252 231 QLP 
Q207 225 253 231 QLN 
D205 225 223 DL     
D206 224 226 DL     
R211 223 221 .26   
R213 222 224 .26   
R2CLP 229 231 .26  
R2CLN 231 230 .26  
R209 253 229 1000   
R210 252 230 1000
*SHARING CIRCUIT
R301 103 3 1.4
R302 203 3 1.4
R303 303 3 1.4
R304 304 3 10
C304 304 5 10E-9
.MODEL DD D(CJO=0.1PF IS=1E-17) 
.MODEL DL D(CJO=3PF IS=1E-13)   
.MODEL QI1 NPN (BF=7.37E-01 IS=8E-16)   
.MODEL QI2 NPN (BF=6.67E-01 IS=8.45E-16)
.MODEL QOP PNP (BF=3.92E+02 IS=1E-14)   
.MODEL QON NPN (BF=3.92E+02 IS=1E-14)   
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
*************
* BEGIN OPAMP MACROMODEL PA75AMP
* REVISION 1 3-MARCH-2004 INITIAL RELEASE
* SYM=PA21
* PINOUT ORDER +IN -IN OUT +V -V
*                1  2   3   4  5
.SUBCKT PA75AMP 1 2 3 4 5 
R4 9 12 7.39E+3 
R3 8 12 7.39E+3 
R1 4 10 8.85E+3 
R2 4 11 8.85E+3 
R5 12 5 111E6   
R6 6 0 100E+3   
R7 7 0 1000     
I2 12 5 16.6E-6 
C1 12 5 2.73E-12
C2 10 11 1E-12  
G1 6 0 11 10 113E-6     
G2 6 0 12 0 6.36E-9     
G3 0 7 0 6 25   
D1 6 0 DD       
D2 0 6 DD       
C3 6 7 4.4E-12  
I1 5 4 10.8E-3  
D3 7 16 DD      
D4 17 7 DD      
V1 18 16 1.63   
V2 17 19 1.63   
I3 4 23 6.3E-3  
I4 24 5 6.3E-3  
Q5 4 23 29 QON  
Q4 4 20 22 QON  
Q6 5 24 30 QOP  
Q3 5 20 21 QOP  
R58 51 20 50    
R8 7 50 50      
C54 20 0 .34E-9 
C4 50 0 .3E-9   
R15 31 3 .76    
E6 18 0 4 0 1   
E7 19 0 5 0 1   
E50 51 0 50 0 1 
Q1 10 1 8 QI1   
Q2 11 2 9 QI2   
Q8 26 28 31 QLP 
Q7 25 27 31 QLN 
D5 25 23 DL     
D6 24 26 DL     
R11 23 21 .26   
R13 22 24 .26   
RCLP 29 31 .26  
RCLN 31 30 .26  
R9 27 29 1000   
R10 28 30 1000
.MODEL DD D(CJO=0.1PF IS=1E-17) 
.MODEL DL D(CJO=3PF IS=1E-13)   
.MODEL QI1 NPN (BF=7.37E-01 IS=8E-16)   
.MODEL QI2 NPN (BF=6.67E-01 IS=8.45E-16)
.MODEL QOP PNP (BF=3.92E+02 IS=1E-14)   
.MODEL QON NPN (BF=3.92E+02 IS=1E-14)   
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
*************
* BEGIN OPAMP MACROMODEL PA75BUF
* REVISION 1 3-MARCH-2004 INITIAL RELEASE
* PINOUT ORDER +IN OUT +V -V
*                1  3   4  5
.SUBCKT PA75BUF 1 3 4 5 
R4 9 12 7.39E+3 
R3 8 12 7.39E+3 
R1 4 10 8.85E+3 
R2 4 11 8.85E+3 
R5 12 5 111E6   
R6 6 0 100E+3   
R7 7 0 1000     
I2 12 5 16.6E-6 
C1 12 5 2.73E-12
C2 10 11 1E-12  
G1 6 0 11 10 113E-6     
G2 6 0 12 0 6.36E-9     
G3 0 7 0 6 25   
D1 6 0 DD       
D2 0 6 DD       
C3 6 7 4.4E-12  
I1 5 4 10.8E-3  
D3 7 16 DD      
D4 17 7 DD      
V1 18 16 1.63   
V2 17 19 1.63   
I3 4 23 6.3E-3  
I4 24 5 6.3E-3  
Q5 4 23 29 QON  
Q4 4 20 22 QON  
Q6 5 24 30 QOP  
Q3 5 20 21 QOP  
R58 51 20 50    
R8 7 50 50      
C54 20 0 .34E-9 
C4 50 0 .3E-9   
R15 31 3 .76    
E6 18 0 4 0 1   
E7 19 0 5 0 1   
E50 51 0 50 0 1 
Q1 10 1 8 QI1   
Q2 11 3 9 QI2   
Q8 26 28 31 QLP 
Q7 25 27 31 QLN 
D5 25 23 DL     
D6 24 26 DL     
R11 23 21 .26   
R13 22 24 .26   
RCLP 29 31 .26  
RCLN 31 30 .26  
R9 27 29 1000   
R10 28 30 1000
.MODEL DD D(CJO=0.1PF IS=1E-17) 
.MODEL DL D(CJO=3PF IS=1E-13)   
.MODEL QI1 NPN (BF=7.37E-01 IS=8E-16)   
.MODEL QI2 NPN (BF=6.67E-01 IS=8.45E-16)
.MODEL QOP PNP (BF=3.92E+02 IS=1E-14)   
.MODEL QON NPN (BF=3.92E+02 IS=1E-14)   
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
*************
* BEGIN OPAMP MACROMODEL PA76
* REVISION 1 15-DECEMBER-2003 INITIAL RELEASE
* SYM=PA21
* PINOUT ORDER +IN -IN OUT +V -V
*                1  2   3   4  5
.SUBCKT PA76 1 2 3 4 5 
R4 9 12 7.39E+3 
R3 8 12 7.39E+3 
R1 4 10 8.85E+3 
R2 4 11 8.85E+3 
R5 12 5 111E6   
R6 6 0 100E+3   
R7 7 0 1000     
I2 12 5 16.6E-6 
C1 12 5 2.73E-12
C2 10 11 1E-12  
G1 6 0 11 10 113E-6     
G2 6 0 12 0 6.36E-9     
G3 0 7 0 6 25   
D1 6 0 DD       
D2 0 6 DD       
C3 6 7 4.4E-12  
I1 5 4 10.8E-3  
D3 7 16 DD      
D4 17 7 DD      
V1 18 16 1.63   
V2 17 19 1.63   
I3 4 23 6.3E-3  
I4 24 5 6.3E-3  
Q5 4 23 29 QON  
Q4 4 20 22 QON  
Q6 5 24 30 QOP  
Q3 5 20 21 QOP  
R58 51 20 50    
R8 7 50 50      
C54 20 0 .34E-9 
C4 50 0 .3E-9   
R15 31 303 .76    
E6 18 0 4 0 1   
E7 19 0 5 0 1   
E50 51 0 50 0 1 
Q1 10 1 8 QI1   
Q2 11 2 9 QI2   
Q8 26 52 31 QLP 
Q7 25 53 31 QLN 
D5 25 23 DL     
D6 24 26 DL     
R11 23 21 .26   
R13 22 24 .26   
RCLP 29 31 .26  
RCLN 31 30 .26  
R9 53 29 1000   
R10 52 30 1000
*BUFFER 1
R104 109 112 7.39E+3 
R103 108 112 7.39E+3 
R101 4 110 8.85E+3 
R102 4 111 8.85E+3 
R105 112 5 111E6   
R106 106 0 100E+3   
R107 107 0 1000     
I102 112 5 16.6E-6 
C101 112 5 2.73E-12
C102 110 111 1E-12  
G101 106 0 111 10 113E-6     
G102 106 0 112 0 6.36E-9     
G103 0 107 0 106 25   
D101 106 0 DD       
D102 0 106 DD       
C103 106 107 4.4E-12  
I101 5 4 10.8E-3  
D103 107 116 DD      
D104 117 107 DD      
V101 118 116 1.63   
V102 117 119 1.63   
I103 4 123 6.3E-3  
I104 124 5 6.3E-3  
Q105 4 123 129 QON  
Q104 4 120 122 QON  
Q106 5 124 130 QOP  
Q103 5 120 121 QOP  
R158 151 120 50    
R108 107 150 50      
C154 120 0 .34E-9 
C104 150 0 .3E-9   
R115 131 103 .76    
E106 118 0 4 0 1   
E107 119 0 5 0 1   
E150 151 0 150 0 1 
Q101 110 303 108 QI1   
Q102 111 103 109 QI2   
Q108 126 152 131 QLP 
Q107 125 153 131 QLN 
D105 125 123 DL     
D106 124 126 DL     
R111 123 121 .26   
R113 122 124 .26   
R1CLP 129 131 .26  
R1CLN 131 130 .26  
R109 153 129 1000   
R110 152 130 1000
*BUFFER2
R204 209 212 7.39E+3 
R203 208 212 7.39E+3 
R201 4 210 8.85E+3 
R202 4 211 8.85E+3 
R205 12 5 111E6   
R206 206 0 100E+3   
R207 207 0 1000     
I202 212 5 16.6E-6 
C201 212 5 2.73E-12
C202 210 211 1E-12  
G201 206 0 211 10 113E-6     
G202 206 0 212 0 6.36E-9     
G203 0 207 0 206 25   
D201 206 0 DD       
D202 0 206 DD       
C203 206 207 4.4E-12  
I201 5 4 10.8E-3  
D203 207 216 DD      
D204 217 207 DD      
V201 218 216 1.63   
V202 217 219 1.63   
I203 4 223 6.3E-3  
I204 224 5 6.3E-3  
Q205 4 223 229 QON  
Q204 4 220 222 QON  
Q206 5 224 230 QOP  
Q203 5 220 221 QOP  
R258 251 220 50    
R208 207 250 50      
C254 220 0 .34E-9 
C204 250 0 .3E-9   
R215 231 203 .76    
E206 218 0 4 0 1   
E207 219 0 5 0 1   
E250 251 0 250 0 1 
Q201 210 303 208 QI1   
Q202 211 203 209 QI2   
Q208 226 252 231 QLP 
Q207 225 253 231 QLN 
D205 225 223 DL     
D206 224 226 DL     
R211 223 221 .26   
R213 222 224 .26   
R2CLP 229 231 .26  
R2CLN 231 230 .26  
R209 253 229 1000   
R210 252 230 1000
*SHARING CIRCUIT
R301 103 3 1.4
R302 203 3 1.4
R303 303 3 1.4
R304 304 3 10
C304 304 5 10E-9
.MODEL DD D(CJO=0.1PF IS=1E-17) 
.MODEL DL D(CJO=3PF IS=1E-13)   
.MODEL QI1 NPN (BF=7.37E-01 IS=8E-16)   
.MODEL QI2 NPN (BF=6.67E-01 IS=8.45E-16)
.MODEL QOP PNP (BF=3.92E+02 IS=1E-14)   
.MODEL QON NPN (BF=3.92E+02 IS=1E-14)   
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
***********
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA21
* BEGIN OPAMP MACROMODEL PA81
* PINOUT ORDER +IN -IN OUT +V -V
*               1   2   3   4  5
.SUBCKT PA81 1 2 3 4 5
J1 10 1 8 JI1
J2 11 2 9 JI2
R3 12 8 4.74E+02
R4 12 9 4.74E+02
I2 12 5 4.40E-04
C1 12 5 2.44E-12
R5 12 5 6.82E+06
R1 4 10 7.24E+02
R2 4 11 7.24E+02
C2 10 11 2.20E-11
I1 4 5 5.11E-03
G1 6 15 11 10 1.38E-03
G2 6 15 12 15 7.77E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 2.20E-11
G3 15 7 15 6 4.07E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 4.70E+00
D4 17 7 DD
V2 17 19 4.70E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 1.16E-10
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 1.19E+01
RCLP 29 31 1.19E+01
RCLN 30 31 1.19E+01
R13 22 24 1.19E+01
D5 23 25 DL
D6 26 24 DL
R9 27 29 1E3
R10 28 30 1E3
I3 18 23 9.47E-04
I4 24 19 9.47E-04
R15 31 3 2.50E+01
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL JI1 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1)
.MODEL JI2 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1.0015)
.MODEL QOP PNP (BF=5.54E+01 IS=1E-14)
.MODEL QON NPN (BF=5.54E+01 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
***********************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA21
* BEGIN OPAMP MACROMODEL PA83
* PINOUT ORDER +IN -IN OUT +V -V
*               1   2   3   4  5
.SUBCKT PA83 1 2 3 4 5
J1 10 1 8 JI1
J2 11 2 9 JI2
R3 12 8 4.74E+02
R4 12 9 4.74E+02
I2 12 5 6.60E-04
C1 12 5 1.57E-12
R5 12 5 4.55E+06
R1 4 10 7.24E+02
R2 4 11 7.24E+02
C2 10 11 2.20E-11
I1 4 5 4.00E-03
G1 6 15 11 10 1.38E-03
G2 6 15 12 15 7.77E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 2.20E-11
G3 15 7 15 6 4.07E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 2.70E+00
D4 17 7 DD
V2 17 19 2.70E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 1.16E-11
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 5.95E+00
RCLP 29 31 5.95E+00
RCLN 30 31 5.95E+00
R13 22 24 5.95E+00
D5 23 25 DL
D6 26 24 DL
R9 27 29 1E3
R10 28 30 1E3
I3 18 23 1.34E-03
I4 24 19 1.34E-03
R15 31 3 4.80E+01
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL JI1 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1)
.MODEL JI2 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1.0015)
.MODEL QOP PNP (BF=7.84E+01 IS=1E-14)
.MODEL QON NPN (BF=7.84E+01 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
********************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA09
* BEGIN OPAMP MACROMODEL PA84
* PINOUT ORDER +IN -IN OUT +V -V COMP COMP
*                1   2  3   4  5   6    7
.SUBCKT PA84 1 2 3 4 5 6 7
* NOTE THAT COMPENSATION DOES NOT CONNECT BETWEEN A COMP PIN
* AND SUPPLY BUT RATHER CONNECTS BETWEEN TWO COMP PINS
* THIS IS A DEVIATION FROM THE PHYSICAL PINOUT OF THE
* REAL PART BUT DOES NOT AFFECT PERFORMANCE OF THE MODEL
J1 10 1 8 JI1
J2 11 2 9 JI2
R3 12 8 5.46E+02
R4 12 9 5.46E+02
I2 12 5 2.00E-03
C1 12 5 1.11E-12
R5 12 5 2.00E+06
R1 4 10 7.96E+02
R2 4 11 7.96E+02
C2 10 11 1.00E-10
I1 4 5 2.55E-03
G1 6 15 11 10 1.26E-03
G2 6 15 12 15 1.26E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 5.00E-12
G3 15 7 15 6 4.48E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 2.20E+00
D4 17 7 DD
V2 17 19 2.20E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 9.20E-11
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 23 29 QON
Q6 5 24 30 QOP
Q7 25 27 31 QLN
Q8 26 28 31 QLP
R11 21 23 1.19E+01
RCLP 29 31 1.19E+01
RCLN 30 31 1.19E+01
R13 22 24 1.19E+01
D5 23 25 DL
D6 26 24 DL
R9 27 29 1E3
R10 28 30 1E3
I3 18 23 9.47E-04
I4 24 19 9.47E-04
R15 31 3 3.75E+01
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL JI1 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1)
.MODEL JI2 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1.0015)
.MODEL QOP PNP (BF=5.54E+01 IS=1E-14)
.MODEL QON NPN (BF=5.54E+01 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
*********************
*REVISION 3 9-SEP-2006
*CORRECTED VOLTAGE SWING AND INCREASED I MAX TO 420MA
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA85
* BEGIN OPAMP MACROMODEL PA85
* PINOUT ORDER +IN -IN CL OUT +V -V COMP COMP
*                1   2  3  33  4  5   6    7
.SUBCKT PA85 1 2 3 33 4 5 6 7
M1 10 1 8 8 MI1
M2 11 2 9 9 MI2
R3 12 8 2.20E+02
R4 12 9 2.20E+02
I2 12 5 7.47E-03
C1 12 5 1.04E-12
R5 12 5 5.35E+06
R1 4 10 3.20E+02
R2 4 11 3.20E+02
C2 10 11 6.22E-11
I1 4 5 1.16E-02
G1 6 15 11 10 3.13E-03
G2 6 15 12 15 9.89E-09
R6 6 15 1.00E+05
D1 6 34 DD
D7 34 15 DD
D2 35 6 DD
D8 15 35 DD
C3 6 7 5.00E-12
G3 15 7 15 6 4.52E-01
R7 7 15 1E3
D3 7 16 DD
V1 18 16 5.9E+00
D4 17 7 DD
V2 17 19 5.9E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 9.36E-12
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 1.89E-03
I4 22 19 1.89E-03
R15 29 3 1.72E+01
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=2.10E-15 RS=1.43E+00)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MI1 NMOS (KP=1.00E-02 IS=3E-16 VTO=1)
.MODEL MI2 NMOS (KP=1.00E-02 IS=3E-16 VTO=0.9990)
.MODEL QOP PNP (BF=2.22E+02 IS=1E-14)
.MODEL QON NPN (BF=2.22E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
******************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA85
* BEGIN OPAMP MACROMODEL PA88
* PINOUT ORDER +IN -IN CL OUT +V -V COMP COMP
*                1   2  3  33  4  5   6    7
.SUBCKT PA88 1 2 3 33 4 5 6 7
M1 10 1 8 8 MI1
M2 11 2 9 9 MI2
R3 12 8 2.95E+03
R4 12 9 2.95E+03
I2 12 5 2.49E-04
C1 12 5 2.86E-13
R5 12 5 3.21E+08
R1 4 10 3.20E+03
R2 4 11 3.20E+03
C2 10 11 3.11E-11
I1 4 5 1.12E-04
G1 6 15 11 10 2.00E-04
G2 6 15 12 15 5.56E-09
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 5.00E-12
G3 15 7 15 6 5.69E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 5.20E+00
D4 17 7 DD
V2 17 19 5.20E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 3.06E-10
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 1.34E-03
I4 22 19 1.34E-03
R15 29 3 5.00E+01
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=1.05E-15 RS=2.86E+00)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MI1 NMOS (KP=4.00E-03 IS=3E-16 VTO=1)
.MODEL MI2 NMOS (KP=4.00E-03 IS=3E-16 VTO=0.9990)
.MODEL QOP PNP (BF=7.84E+01 IS=1E-14)
.MODEL QON NPN (BF=7.84E+01 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
*********************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA85
* BEGIN OPAMP MACROMODEL PA89
* PINOUT ORDER +IN -IN CL OUT +V -V COMP COMP
*                1   2  3  33  4  5   6    7
.SUBCKT PA89 1 2 3 33 4 5 6 7
M1 10 1 8 8 MI1
M2 11 2 9 9 MI2
R3 12 8 2.48E+02
R4 12 9 2.48E+02
I2 12 5 3.20E-04
C1 12 5 1.33E-12
R5 12 5 3.75E+07
R1 4 10 4.98E+02
R2 4 11 4.98E+02
C2 10 11 1.07E-10
I1 4 5 3.32E-03
G1 6 15 11 10 2.01E-03
G2 6 15 12 15 3.19E-08
R6 6 15 1.00E+05
D1 6 34 DD
D7 34 15 DD
D2 35 6 DD
D8 15 35 DD
C3 6 7 5.00E-12
G3 15 7 15 6 1.25E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 1.12E+01
D4 17 7 DD
V2 17 19 1.12E+01
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 1.15E-10
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 1.16E-03
I4 22 19 1.16E-03
R15 29 3 6.00E+01
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=7.88E-16 RS=3.81E+00)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MI1 NMOS (KP=4.00E-03 IS=3E-16 VTO=1)
.MODEL MI2 NMOS (KP=4.00E-03 IS=3E-16 VTO=0.9990)
.MODEL QOP PNP (BF=6.79E+01 IS=1E-14)
.MODEL QON NPN (BF=6.79E+01 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
******************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA85
* BEGIN OPAMP MACROMODEL PA90
* NOTE THAT IQ PIN IS NOT MODELED
* PINOUT ORDER +IN -IN CL OUT +V -V COMP COMP
*                1   2  3  33  4  5   6    7
.SUBCKT PA90 1 2 3 33 4 5 6 7
J1 10 1 8 JI1
J2 11 36 9 JI2
R3 12 8 8.88E+01
R4 12 9 8.88E+01
I2 12 5 1.62E-03
C1 12 5 4.75E-14
R5 12 5 3.08E+06
R1 4 10 3.39E+02
R2 4 11 3.39E+02
C2 10 11 5.88E-11
I1 4 5 5.80E-03
G1 6 15 11 10 2.95E-03
G2 37 15 12 15 1.00E-04
LCM 37 38 1.0E-06
RCM 15 38 1.0
ECA 2 36 37 15 1.0
R6 6 15 7.51E+04
D1 6 34 DD
D7 34 15 DD
D2 35 6 DD
D8 15 35 DD
C3 6 7 4.70E-12
G3 15 7 15 6 2.85E-01
R7 7 15 1E3
D3 7 16 DD
V1 18 16 4.20E+00
D4 17 7 DD
V2 17 19 4.20E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 5.60E-12
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 2.58E-03
I4 22 19 2.58E-03
R15 29 3 8.67E+00
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=3.88E-15 RS=7.72E-01)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL JI1 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1 KF=7.0E-18)
.MODEL JI2 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1.0020 KF=7.0E-18)
.MODEL QOP PNP (BF=1.51E+02 IS=1E-14)
.MODEL QON NPN (BF=1.51E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
******************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA85
* BEGIN OPAMP MACROMODEL PA91
* NOTE THAT IQ PIN IS NOT MODELED
* PINOUT ORDER +IN -IN CL OUT +V -V COMP COMP
*                1   2  3  33  4  5   6    7
.SUBCKT PA91 1 2 3 33 4 5 6 7
J1 10 1 8 JI1
J2 11 36 9 JI2
R3 12 8 8.88E+01
R4 12 9 8.88E+01
I2 12 5 1.62E-03
C1 12 5 4.75E-14
R5 12 5 3.08E+06
R1 4 10 3.39E+02
R2 4 11 3.39E+02
C2 10 11 5.88E-11
I1 4 5 5.80E-03
G1 6 15 11 10 2.95E-03
G2 37 15 12 15 1.00E-04
LCM 37 38 1.0E-06
RCM 15 38 1.0
ECA 2 36 37 15 1.0
R6 6 15 7.51E+04
D1 6 34 DD
D7 34 15 DD
D2 35 6 DD
D8 15 35 DD
C3 6 7 4.70E-12
G3 15 7 15 6 2.85E-01
R7 7 15 1E3
D3 7 16 DD
V1 18 16 4.20E+00
D4 17 7 DD
V2 17 19 4.20E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 5.60E-12
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 2.58E-03
I4 22 19 2.58E-03
R15 29 3 8.67E+00
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=3.88E-15 RS=7.72E-01)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL JI1 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1 KF=7.0E-18)
.MODEL JI2 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1.0020 KF=7.0E-18)
.MODEL QOP PNP (BF=1.51E+02 IS=1E-14)
.MODEL QON NPN (BF=1.51E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
******************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA85
* BEGIN OPAMP MACROMODEL PA92
* NOTE THAT IQ PIN IS NOT MODELED
* PINOUT ORDER +IN -IN CL OUT +V -V COMP COMP
*                1   2  3  33  4  5   6    7
.SUBCKT PA92 1 2 3 33 4 5 6 7
J1 10 1 8 JI1
J2 11 36 9 JI2
R3 12 8 5.17E+02
R4 12 9 5.17E+02
I2 12 5 7.20E-04
C1 12 5 4.32E-13
R5 12 5 9.72E+07
C7 9 41 1.71E-10
RZ1 12 40 5.17E+01
C8 8 40 1.71E-10
RZ2 12 41 5.17E+01
R1 4 10 5.42E+02
R2 4 11 5.42E+02
C2 10 11 3.68E-11
I1 4 5 -2.86E-03
G1 6 15 11 10 1.85E-03
G2 37 15 12 15 1.00E-04
LCM 37 38 1.0E-06
RCM 15 38 1.0
ECA 2 36 37 15 1.0
R6 6 15 1.00E+05
D1 6 34 DD
D7 34 15 DD
D2 35 6 DD
D8 15 35 DD
C3 6 7 4.70E-12
G3 15 7 15 6 3.42E-01
R7 7 15 1E3
D3 7 16 DD
V1 18 16 7.10E+00
D4 17 7 DD
V2 17 19 7.10E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 42 50
C4 42 15 2.80E-11
R11 20 42 50
C5 20 15 4.55E-10
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 333
R10 28 3 333
I3 18 21 1.23E-02
I4 22 19 1.23E-02
R15 29 3 5.43E-01
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=8.92E-14 RS=3.36E-02)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL JI1 NJF (BETA=4.00E-02 IS=3E-16 VTO=-1 KF=7.0E-18)
.MODEL JI2 NJF (BETA=4.00E-02 IS=3E-16 VTO=-1.0020 KF=7.0E-18)
.MODEL QOP PNP (BF=7.23E+02 IS=1E-14)
.MODEL QON NPN (BF=7.23E+02 IS=1E-14)
.MODEL QLN NPN (BF=200 IS=6E-13)
.MODEL QLP PNP (BF=200 IS=6E-13)
* END OF OPAMP MACROMODEL
.ENDS
******************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA85
* BEGIN OPAMP MACROMODEL PA93
* NOTE THAT IQ PIN IS NOT MODELED
* PINOUT ORDER +IN -IN CL OUT +V -V COMP COMP
*                1   2  3  33  4  5   6    7
.SUBCKT PA93 1 2 3 33 4 5 6 7
J1 10 1 8 JI1
J2 11 36 9 JI2
R3 12 8 5.17E+02
R4 12 9 5.17E+02
I2 12 5 7.20E-04
C1 12 5 4.32E-13
R5 12 5 9.72E+07
C7 9 41 3.08E-10
RZ1 12 40 5.17E+01
C8 8 40 3.08E-10
RZ2 12 41 5.17E+01
R1 4 10 5.42E+02
R2 4 11 5.42E+02
C2 10 11 5.88E-11
I1 4 5 -6.91E-03
G1 6 15 11 10 1.85E-03
G2 37 15 12 15 1.00E-04
LCM 37 38 1.0E-06
RCM 15 38 1.0
ECA 2 36 37 15 1.0
R6 6 15 1.00E+05
D1 6 34 DD
D7 34 15 DD
D2 35 6 DD
D8 15 35 DD
C3 6 7 4.70E-12
G3 15 7 15 6 3.42E-01
R7 7 15 1E3
D3 7 16 DD
V1 18 16 6.20E+00
D4 17 7 DD
V2 17 19 6.20E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 42 50
C4 42 15 2.80E-11
R11 20 42 50
C5 20 15 6.37E-10
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 333
R10 28 3 333
I3 18 21 1.64E-02
I4 22 19 1.64E-02
R15 29 3 3.43E-01
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=1.57E-13 RS=1.90E-02)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL JI1 NJF (BETA=4.00E-02 IS=3E-16 VTO=-1 KF=7.0E-18)
.MODEL JI2 NJF (BETA=4.00E-02 IS=3E-16 VTO=-1.0020 KF=7.0E-18)
.MODEL QOP PNP (BF=9.60E+02 IS=1E-14)
.MODEL QON NPN (BF=9.60E+02 IS=1E-14)
.MODEL QLN NPN (BF=200 IS=6E-13)
.MODEL QLP PNP (BF=200 IS=6E-13)
* END OF OPAMP MACROMODEL
.ENDS
******************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA85
* BEGIN OPAMP MACROMODEL PA94
* PINOUT ORDER +IN -IN CL OUT +V -V COMP COMP
*                1   2  3  33  4  5   6    7
.SUBCKT PA94 1 2 3 33 4 5 6 7
J1 10 1 8 JI1
J2 11 2 9 JI2
R3 12 8 5.07E+01
R4 12 9 5.07E+01
I2 12 5 4.10E-03
C1 12 5 5.49E-14
R5 12 5 3.24E+07
R1 4 10 1.22E+02
R2 4 11 1.22E+02
C2 10 11 1.87E-10
I1 4 5 1.23E-02
G1 6 15 11 10 8.20E-03
G2 6 15 12 15 1.03E-07
R6 6 15 1.00E+05
D1 6 34 DD
D7 34 15 DD
D2 35 6 DD
D8 15 35 DD
C3 6 7 3.24E-12
G3 15 7 15 6 6.86E-01
R7 7 15 1E3
D3 7 16 DD
V1 18 16 8.20E+00
D4 17 7 DD
V2 17 19 8.20E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 2.23E-10
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 1.89E-03
I4 22 19 1.89E-03
R15 29 3 1.50E+02
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=2.10E-15 RS=1.43E+00)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL JI1 NJF (BETA=1.40E-02 IS=3E-16 VTO=-1)
.MODEL JI2 NJF (BETA=1.40E-02 IS=3E-16 VTO=-1.0050)
.MODEL QOP PNP (BF=1.11E+02 IS=1E-14)
.MODEL QON NPN (BF=1.11E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
******************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA85
* BEGIN OPAMP MACROMODEL PA95
* PINOUT ORDER +IN -IN CL OUT +V -V COMP COMP
*                1   2  3  33  4  5   6    7
.SUBCKT PA95 1 2 3 33 4 5 6 7
J1 10 1 8 JI1
J2 11 36 9 JI2
R3 12 8 9.78E+02
R4 12 9 9.78E+02
I2 12 5 2.40E-04
C1 12 5 8.02E-14
R5 12 5 5.40E+08
C7 9 41 1.63E-12
RZ1 12 40 9.78E+01
C8 8 40 1.63E-12
RZ2 12 41 9.78E+01
R1 4 10 1.00E+03
R2 4 11 1.00E+03
C2 10 11 1.13E-11
I1 4 5 -4.60E-04
G1 6 15 11 10 9.97E-04
G2 37 15 12 15 1.26E-05
LCM 37 38 1.0E-06
RCM 15 38 1.0
ECA 2 36 37 15 1.0
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 3.24E-12
G3 15 7 15 6 7.97E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 9.20E+00
D4 17 7 DD
V2 17 19 9.20E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 42 50
C4 42 15 2.81E-11
R11 20 42 50
C5 20 15 4.55E-10
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 333
R10 28 3 333
I3 18 21 1.89E-03
I4 22 19 1.89E-03
R15 29 3 1.44E+02
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=2.10E-15 RS=1.43E+00)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL JI1 NJF (BETA=4.00E-02 IS=3E-16 VTO=-1 KF=7.0E-18)
.MODEL JI2 NJF (BETA=4.00E-02 IS=3E-16 VTO=-1.0005 KF=7.0E-18)
.MODEL QOP PNP (BF=1.11E+02 IS=1E-14)
.MODEL QON NPN (BF=1.11E+02 IS=1E-14)
.MODEL QLN NPN (BF=200 IS=6E-13)
.MODEL QLP PNP (BF=200 IS=6E-13)
* END OF OPAMP MACROMODEL
.ENDS
******************
* REVISION 1 FEB 15 2007 INITIAL RELEASE
* SYMPOL PA85
* BEGIN MODEL PA96
* PINOUT ORDER +IN -IN CL OUT +V -V COMP COMP
* PINOUT ORDER  4   5   2  1   3  6   7    8
* NOTE THAT THIS MODEL DOES NOT PERFORM THE
* BANDWIDTH FALLOFF AT LOWER +SUPPLY VOLTAGE
* AS SHOWN IN THE DATA SHEET
.SUBCKT PA96 4 5 2 1 3 6 7 8
R83 9 10 10
R85 11 12 10
R86 7 13 100
R93 6 14 311
R94 6 15 129
D6 13 16 N5242
E2 17 18 3 6 -2.66E-3
D8 19 0 DD
I1 0 19 1E-3
V16 19 20 0.7
E3 21 0 20 0 -571
R98 0 20 1E6
R99 0 21 1E6
E4 8 9 22 0 2.5E-3
E5 18 11 22 0 -2.5E-3
V17 21 22 27
R100 0 22 1E6
D9 17 8 DZ
J2 23 5 24 N912
J3 13 25 26 N912
R101 27 24 43
R102 27 26 43
Q13 23 28 29 Q907C
Q14 13 23 30 Q907C
R103 29 16 115
R104 30 16 115
V18 25 31 -3E-3
R109 32 16 39
Q15 33 2 1 Q222
Q16 18 2 1 Q908
E99 34 35 36 0 0.01
R118 36 37 1E6
R119 0 36 100
C25 37 36 1E-12
E100 37 0 3 0 1
R120 35 34 1E9
E101 35 38 39 0 -0.01
R121 39 40 1E6
R122 0 39 100
C26 40 39 20E-12
E102 40 0 6 0 1
R123 38 35 1E9
E103 38 41 42 0 -0.125
R124 42 43 1E6
R125 0 42 100
C27 43 42 20E-12
E104 43 0 44 0 1
R126 41 38 1E9
E105 41 4 45 46 4
D17 45 0 DVN
I7 0 45 100E-6
D18 46 0 DVN
I8 0 46 100E-6
R127 4 41 1E9
E106 47 0 34 0 1
E107 48 0 5 0 1
R128 44 47 1E3
R129 44 48 1E3
R130 6 3 12E6
E108 31 34 22 0 31E-6
R131 34 31 1E9
C28 5 0 4E-12
C29 34 0 4E-12
I9 3 6 2.3E-3
R133 18 17 1E9
X10 18 6 15 D3545
X11 49 14 50 D3545
X12 51 13 32 P2450
R145 52 2 0.006
R148 53 2 0.031
C31 8 18 10E-9
C32 7 8 1E-12
M1 6 12 53 53 VP0335 L=2.5E-6 W=8.85E-2
M2 3 10 52 52 VN0335 L=3.0E-6 W=8.12E-2
Q17 50 54 14 Q222
D21 6 54 DZ1
I10 3 54 0.5E-3
X13 51 33 8 D3545
R149 8 33 420
C34 23 13 10E-12
R151 28 23 200
V27 27 49 0
V28 3 16 0
.MODEL DZ1 D(IS=5E-11 RS=14 BV=2.81 IBV=6E-4 KF=1E-15)
.MODEL DVN D KF=5E-16
.MODEL DD D
.MODEL Q222 NPN IS=2E-13
.MODEL Q908 PNP IS=1E-13
.MODEL DZ D BV=6.043 IBV=0.001 RS=5
.MODEL N912 NJF VTO=-3 BETA=3.2E-3 RS=12 RD=50
+ IS=1E-18 LAMBDA=3E-4 CGS=10E-12 CGD=0.5E-12
.MODEL N5242 D IS=1E-15 RS=5 N=1 BV=12 IBV=1E-4
.MODEL Q907C PNP IS=1.1E-13 BF=150 BR=6 NF=1.2
+ RC=1 IKF=0.1 VAF=340 XTB=1.5 NE=1.8 ISE=1.5E-13
+ CJE=20E-12 VJE=0.8 MJE=1.2 CJC=15E-12 VJC=0.57
+ MJC=0.3 TF=0.5E-9 TR=35E-9
.MODEL VN0335 NMOS (LEVEL=3 RS=0.11 NSUB=5.0E15
+DELTA=0.1 KAPPA=0.10123 TPG=1  CGDO=1.2E-10
+RD=7.0 VTO=3.00   VMAX=1.0E7  ETA=0.0223089
+NFS=6.6E10 TOX=1.0E-7 LD=1.698E-9 UO=862.425
+XJ=6.4666E-7 THETA=1.0E-5 CGSO=2.1E-9
+CBD=40E-12)
.MODEL VP0335 PMOS (LEVEL=3 RS=0.25 NSUB=5.0E15
+DELTA=0.1 KAPPA=0.10123 TPG=-1 CGDO=1.2E-10
+RD=8.2 VTO=-3.00 VMAX=1.0E7 ETA=0.0223089
+NFS=6.6E10 TOX=1.0E-7 LD=1.698E-9 UO=862.425
+XJ=6.4666E-7 THETA=1.0E-5 CGSO=2.1E-9
+CBD=40E-12)
.ENDS PA96
.SUBCKT D3545 10 20 30
M1 10 20 30 30 DMOS L=1U W=1U
CGS 20 30 43E-12
.MODEL DMOS NMOS LEVEL=3 VMAX=9E5 THETA=6E-3
+ ETA=2E-4 VTO=-1.53 KP=0.07 RS=2 RD=19)
.ENDS
.SUBCKT P2450 10 20 30
M1 10 20 30 30 DMOS L=1U W=1U
RDS 10 30 1E6
CGS 20 30 100E-12
CDG 10 20 1E-12
.MODEL DMOS PMOS LEVEL=3 VMAX=9E5 THETA=60E-3
+ ETA=2E-3 VTO=-2 KP=0.07 RS=3 RD=10)
.ENDS
* END MODEL PA96
************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA09
* BEGIN OPAMP MACROMODEL PA97
* PINOUT ORDER +IN -IN OUT +V -V COMP COMP
*                1   2  3   4  5   6    7
.SUBCKT PA97 1 2 3 4 5 6 7
J1 10 1 8 JI1
J2 11 2 9 JI2
R3 12 8 7.05E+02
R4 12 9 7.05E+02
I2 12 5 1.06E-04
C1 12 5 1.34E-13
R5 12 5 1.24E+09
R1 4 10 9.55E+02
R2 4 11 9.55E+02
C2 10 11 8.34E-11
I1 5 4 4.64E-05
RI1 4 5 8.90E6
G1 6 15 11 10 1.05E-03
G2 6 15 12 15 1.32E-08
R6 6 15 1.00E+05
D1 6 15 DD
D2 15 6 DD
C3 6 7 3.24E-12
G3 15 7 15 6 9.55E+00
R7 7 15 1E3
D3 7 16 DD
V1 18 16 1.40E+01
D4 17 7 DD
V2 17 19 1.02E+01
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 9.44E-10
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
I3 18 21 5.19E-04
I4 22 19 5.19E-04
R15 29 3 9.09E+01
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=1.57E-16 RS=1.90E+01)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL JI1 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1)
.MODEL JI2 NJF (BETA=4.00E-03 IS=3E-16 VTO=-1.0005)
.MODEL QOP PNP (BF=3.04E+01 IS=1E-14)
.MODEL QON NPN (BF=3.04E+01 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
******************
*REVISION 2 18-MAR-2002
*REDUCED INTERACTION OF SLEW RATE WITH CHANGING SUPPLY.
*SYM=PA85
* BEGIN OPAMP MACROMODEL PA98
* PINOUT ORDER +IN -IN CL OUT +V -V COMP COMP
*                1   2  3  33  4  5   6    7
.SUBCKT PA98 1 2 3 33 4 5 6 7
M1 10 1 8 8 MI1
M2 11 2 9 9 MI2
R3 12 8 2.20E+02
R4 12 9 2.20E+02
I2 12 5 7.47E-03
C1 12 5 1.04E-12
R5 12 5 5.35E+06
R1 4 10 3.20E+02
R2 4 11 3.20E+02
C2 10 11 6.22E-11
I1 4 5 1.06E-02
G1 6 15 11 10 3.13E-03
G2 6 15 12 15 9.89E-09
R6 6 15 1.00E+05
D1 6 34 DD
D7 34 15 DD
D2 35 6 DD
D8 15 35 DD
C3 6 7 5.00E-12
G3 15 7 15 6 4.52E-01
R7 7 15 1E3
D3 7 16 DD
V1 18 16 8.70E+00
D4 17 7 DD
V2 17 19 8.70E+00
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
R8 7 20 50
C4 20 15 9.36E-12
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 1.89E-03
I4 22 19 1.89E-03
R15 29 3 2.22E+01
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=10PF IS=2.10E-15 RS=1.43E+00)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MI1 NMOS (KP=1.00E-02 IS=3E-16 VTO=1)
.MODEL MI2 NMOS (KP=1.00E-02 IS=3E-16 VTO=0.9950)
.MODEL QOP PNP (BF=1.11E+02 IS=1E-14)
.MODEL QON NPN (BF=1.11E+02 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-14)
.MODEL QLP PNP (BF=100 IS=1E-14)
* END OF OPAMP MACROMODEL
.ENDS
**********************
*SYM=PB50
* BEGIN OPAMP MACROMODEL PB50
* PINOUT ORDER  IN COM CL OUT +V -V GAIN COMP
*                1   2  3  33  4  5  11   10
.SUBCKT PB50 1 2 3 33 4 5 11 10
Q1 8 1 10 QIN
Q2 8 9 4 QIP
I1 10 5 1.4E-3
RZ1 10 5 200E3
I2 7 5 5E-3
I9 4 5 8E-3
RI9 4 5 25E3
R1 1 2 50E3
R2 2 10 3100
R3 10 11 6200
M1 7 8 13 13 MSS
RG2 13 4 300
CE1 13 4 220E-12
R4 7 5 200E3
C1 7 0 53E-12
R5 4 9 332
R6 8 9 4400
D3 7 16 DD
V1 18 16 5.7
D4 17 7 DD
V2 17 19 5.7
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
E9 12 0 7 0 1
R8 12 20 50
C4 20 15 530E-12
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 2.5E-03
I4 22 19 2.5E-03
R15 29 3 2.25
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=30PF IS=2.10E-14 RS=1.43E-01)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MSS PMOS (KP=1E-02 IS=3E-16 VTO=-2.5)
.MODEL QOP PNP (BF=1200 IS=1E-14)
.MODEL QON NPN (BF=1200 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-11)
.MODEL QLP PNP (BF=100 IS=1E-11)
.MODEL QIN NPN (BF=100 IS=4E-16)
.MODEL QIP PNP (BF=100 IS=4E-16)
* END OF OPAMP MACROMODEL
.ENDS
******************
*SYM=PB50
* BEGIN OPAMP MACROMODEL PB51
* PINOUT ORDER  IN COM CL OUT +V -V GAIN COMP
*                1   2  3  33  4  5  11   10
.SUBCKT PB51 1 2 3 33 4 5 11 10
Q1 8 1 10 QIN
Q2 8 9 4 QIP
I1 10 5 1.4E-3
RZ1 10 5 200E3
I2 7 5 5E-3
I9 4 5 8E-3
RI9 4 5 25E3
R1 1 2 50E3
R2 2 10 3100
R3 10 11 6200
M1 7 8 13 13 MSS
RG2 13 4 300
CE1 13 4 220E-12
R4 7 5 200E3
C1 7 0 53E-12
R5 4 9 332
R6 8 9 4400
D3 7 16 DD
V1 18 16 5.7
D4 17 7 DD
V2 17 19 5.7
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
E9 12 0 7 0 1
R8 12 20 50
C4 20 15 530E-12
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 2.5E-03
I4 22 19 2.5E-03
R15 29 3 2.25
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=30PF IS=2.10E-14 RS=1.43E-01)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MSS PMOS (KP=1E-02 IS=3E-16 VTO=-2.5)
.MODEL QOP PNP (BF=700 IS=1E-14)
.MODEL QON NPN (BF=700 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-11)
.MODEL QLP PNP (BF=100 IS=1E-11)
.MODEL QIN NPN (BF=100 IS=4E-16)
.MODEL QIP PNP (BF=100 IS=4E-16)
* END OF OPAMP MACROMODEL
.ENDS
********************
*SYM=PB50
* BEGIN OPAMP MACROMODEL PB51A
* PINOUT ORDER  IN COM CL OUT +V -V GAIN COMP
*                1   2  3  33  4  5  11   10
.SUBCKT PB51A 1 2 3 33 4 5 11 10
Q1 8 1 10 QIN
Q2 8 9 4 QIP
I1 10 5 1.4E-3
RZ1 10 5 200E3
I2 7 5 5E-3
I9 4 5 8E-3
RI9 4 5 25E3
R1 1 2 50E3
R2 2 10 3100
R3 10 11 6200
M1 7 8 13 13 MSS
RG2 13 4 300
CE1 13 4 220E-12
R4 7 5 200E3
C1 7 0 36E-12
R5 4 9 332
R6 8 9 4400
D3 7 16 DD
V1 18 16 5.7
D4 17 7 DD
V2 17 19 5.7
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
E9 12 0 7 0 1
R8 12 20 50
C4 20 15 355E-12
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 2.5E-03
I4 22 19 2.5E-03
R15 29 3 2.25
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=30PF IS=2.10E-14 RS=1.43E-01)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MSS PMOS (KP=1E-02 IS=3E-16 VTO=-2.5)
.MODEL QOP PNP (BF=933 IS=1E-14)
.MODEL QON NPN (BF=933 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-11)
.MODEL QLP PNP (BF=100 IS=1E-11)
.MODEL QIN NPN (BF=100 IS=4E-16)
.MODEL QIP PNP (BF=100 IS=4E-16)
* END OF OPAMP MACROMODEL
.ENDS
******************
*SYM=PB50
* BEGIN OPAMP MACROMODEL PB58
* PINOUT ORDER  IN COM CL OUT +V -V GAIN COMP
*                1   2  3  33  4  5  11   10
.SUBCKT PB58 1 2 3 33 4 5 11 10
Q1 8 1 10 QIN
Q2 8 9 4 QIP
I1 10 5 1.4E-3
RZ1 10 5 200E3
I2 7 5 5E-3
I9 4 5 8E-3
RI9 4 5 25E3
R1 1 2 50E3
R2 2 10 3100
R3 10 11 6200
M1 7 8 13 13 MSS
RG2 13 4 300
CE1 13 4 220E-12
R4 7 5 200E3
C1 7 0 53E-12
R5 4 9 332
R6 8 9 4400
D3 7 16 DD
V1 18 16 5.7
D4 17 7 DD
V2 17 19 5.7
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
E9 12 0 7 0 1
R8 12 20 50
C4 20 15 530E-12
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 2.5E-03
I4 22 19 2.5E-03
R15 29 3 2.25
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=30PF IS=2.10E-14 RS=1.43E-01)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MSS PMOS (KP=1E-02 IS=3E-16 VTO=-2.5)
.MODEL QOP PNP (BF=700 IS=1E-14)
.MODEL QON NPN (BF=700 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-11)
.MODEL QLP PNP (BF=100 IS=1E-11)
.MODEL QIN NPN (BF=100 IS=4E-16)
.MODEL QIP PNP (BF=100 IS=4E-16)
* END OF OPAMP MACROMODEL
.ENDS
********************
*SYM=PB50
* BEGIN OPAMP MACROMODEL PB58A
* PINOUT ORDER  IN COM CL OUT +V -V GAIN COMP
*                1   2  3  33  4  5  11   10
.SUBCKT PB58A 1 2 3 33 4 5 11 10
Q1 8 1 10 QIN
Q2 8 9 4 QIP
I1 10 5 1.4E-3
RZ1 10 5 200E3
I2 7 5 5E-3
I9 4 5 8E-3
RI9 4 5 25E3
R1 1 2 50E3
R2 2 10 3100
R3 10 11 6200
M1 7 8 13 13 MSS
RG2 13 4 300
CE1 13 4 220E-12
R4 7 5 200E3
C1 7 0 36E-12
R5 4 9 332
R6 8 9 4400
D3 7 16 DD
V1 18 16 5.7
D4 17 7 DD
V2 17 19 5.7
RE1 15 0 0.001
E2 18 0 4 0 1
E3 19 0 5 0 1
E9 12 0 7 0 1
R8 12 20 50
C4 20 15 355E-12
Q3 19 20 21 QOP
Q4 18 20 22 QON
Q5 4 21 29 QON
Q6 5 22 29 QOP
Q7 25 27 33 QLN
Q8 26 28 33 QLP
D5 21 25 DL
D6 26 22 DL
R9 27 3 1E3
R10 28 3 1E3
I3 18 21 2.5E-03
I4 22 19 2.5E-03
R15 29 3 2.25
DC1 29 4 DO
DC2 5 29 DO
.MODEL DO D(CJO=30PF IS=2.10E-14 RS=1.43E-01)
.MODEL DD D(CJO=0.1PF IS=1E-17)
.MODEL DL D(CJO=3PF IS=1E-13)
.MODEL MSS PMOS (KP=1E-02 IS=3E-16 VTO=-2.5)
.MODEL QOP PNP (BF=933 IS=1E-14)
.MODEL QON NPN (BF=933 IS=1E-14)
.MODEL QLN NPN (BF=100 IS=1E-11)
.MODEL QLP PNP (BF=100 IS=1E-11)
.MODEL QIN NPN (BF=100 IS=4E-16)
.MODEL QIP PNP (BF=100 IS=4E-16)
* END OF OPAMP MACROMODEL
.ENDS
**********************
